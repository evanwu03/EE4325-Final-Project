/home/010/e/eb/ebw220000/cad/EE4325_UART_Project/gf65/gf65.lef