* File: OAI22.pex.sp
* Created: Sun May 11 15:40:51 2025
* Program "Calibre xRC"
* Version "v2024.4_12.9"
* 
.include "OAI22.pex.sp.pex"
.subckt OAI22  OUT VSS VDD A B D C
* 
* C	C
* D	D
* B	B
* A	A
* VDD	VDD
* VSS	VSS
* OUT	OUT
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=9.34934e-12
+ PERIM=1.2258e-05
XMMN1 N_OUT_MMN1_d N_A_MMN1_g N_NET3_MMN1_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.3944e-13 AS=9.296e-14 PD=1.058e-06 PS=1.452e-06 NRD=0.183333
+ NRS=0.182143 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.66e-07
+ SB=2.019e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN0 N_OUT_MMN1_d N_B_MMN0_g N_NET3_MMN0_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.3944e-13 AS=1.2768e-13 PD=1.058e-06 PS=1.016e-06 NRD=0.705952
+ NRS=0.390476 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=7.29e-07
+ SB=1.456e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN3 N_NET3_MMN0_s N_D_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2768e-13 AS=1.6296e-13 PD=1.016e-06 PS=1.142e-06 NRD=0.42381
+ NRS=0.502976 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.25e-06
+ SB=9.35e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN2 N_NET3_MMN2_d N_C_MMN2_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.6128e-13 AS=1.6296e-13 PD=1.696e-06 PS=1.142e-06 NRD=0.181548
+ NRS=0.53631 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.897e-06
+ SB=2.88e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMP0 NET2 N_A_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.37795e-13 AS=1.5853e-13 PD=1.453e-06 PS=2.242e-06 NRD=0.260733
+ NRS=0.104712 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.66e-07
+ SB=2.019e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=3.5335e-14
+ PANW6=2.674e-14 PANW7=0 PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP2 N_OUT_MMP2_d N_B_MMP2_g NET2 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.1774e-13 AS=2.37795e-13 PD=1.411e-06 PS=1.453e-06 NRD=0.239791
+ NRS=0.260733 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=7.29e-07
+ SB=1.456e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=9.0935e-14 PANW10=1.3442e-13
XMMP3 N_OUT_MMP2_d N_D_MMP3_g NET1 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.1774e-13 AS=2.77905e-13 PD=1.411e-06 PS=1.537e-06 NRD=0.237696
+ NRS=0.304712 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.25e-06
+ SB=9.35e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=9.0935e-14 PANW10=1.3442e-13
XMMP1 NET1 N_C_MMP1_g N_VDD_MMP1_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.77905e-13 AS=2.7504e-13 PD=1.537e-06 PS=2.486e-06 NRD=0.304712
+ NRS=0.197906 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.897e-06
+ SB=2.88e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=6.2075e-14 PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
*
.include "OAI22.pex.sp.OAI22.pxi"
*
.ends
*
*
