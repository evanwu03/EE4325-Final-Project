* File: DFF.pex.sp
* Created: Thu May  8 20:09:47 2025
* Program "Calibre xRC"
* Version "v2024.4_12.9"
* 
.include "DFF.pex.sp.pex"
.subckt DFF  VSS Q VDD CLK R D
* 
* D	D
* R	R
* CLK	CLK
* VDD	VDD
* Q	Q
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=2.71981e-11
+ PERIM=2.3178e-05
XMMN2 N_CLK-_MMN2_d N_CLK_MMN2_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.6e-07 AD=9.632e-14 AS=1.2572e-13 PD=1.464e-06 PS=1.009e-06
+ NRD=0.185714 NRS=0.601786 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.72e-07 SB=6.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN1 N_CLK+_MMN1_d N_CLK-_MMN1_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.6e-07 AD=9.464e-14 AS=1.2572e-13 PD=1.458e-06 PS=1.009e-06
+ NRD=0.183929 NRS=0.2 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=6.86e-07
+ SB=1.69e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN5 N_B_MMN5_d N_R_MMN5_g N_VSS_MMN5_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.3944e-13 AS=9.296e-14 PD=1.058e-06 PS=1.452e-06 NRD=0.375
+ NRS=0.183929 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.66e-07
+ SB=5e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0
+ PANW9=8.385e-15 PANW10=2.8015e-14
XMMN4 N_B_MMN5_d N_A_MMN4_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.3944e-13 AS=1.274e-13 PD=1.058e-06 PS=1.015e-06 NRD=0.514286
+ NRS=0.226786 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=7.29e-07
+ SB=5e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0
+ PANW9=8.385e-15 PANW10=2.8015e-14
XMMN0 NET1 N_D_MMN0_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.3636e-13 AS=1.274e-13 PD=1.047e-06 PS=1.015e-06 NRD=0.434821
+ NRS=0.585714 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.249e-06
+ SB=4.651e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN3 N_A_MMN3_d N_CLK-_MMN3_g NET1 N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2796e-13 AS=1.3636e-13 PD=1.017e-06 PS=1.047e-06 NRD=0.407143
+ NRS=0.434821 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.801e-06
+ SB=4.099e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN7 N_A_MMN3_d N_CLK+_MMN7_g NET2 N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2796e-13 AS=1.2824e-13 PD=1.017e-06 PS=1.018e-06 NRD=0.408929
+ NRS=0.408929 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.323e-06
+ SB=3.577e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN6 NET2 N_B_MMN6_g N_VSS_MMN6_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2824e-13 AS=1.274e-13 PD=1.018e-06 PS=1.015e-06 NRD=0.408929
+ NRS=0.467857 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.846e-06
+ SB=3.054e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN8 NET3 N_B_MMN8_g N_VSS_MMN6_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.274e-13 AS=1.274e-13 PD=1.015e-06 PS=1.015e-06 NRD=0.40625
+ NRS=0.344643 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.366e-06
+ SB=2.534e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN9 N_C_MMN9_d N_CLK+_MMN9_g NET3 N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2768e-13 AS=1.274e-13 PD=1.016e-06 PS=1.015e-06 NRD=0.433929
+ NRS=0.40625 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.886e-06
+ SB=2.014e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN13 N_C_MMN9_d N_CLK-_MMN13_g NET4 N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2768e-13 AS=6.328e-14 PD=1.016e-06 PS=7.86e-07 NRD=0.380357
+ NRS=0.201786 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=4.407e-06
+ SB=1.493e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN12 NET4 N_E_MMN12_g N_VSS_MMN12_s N_VSS_D0_noxref_pos NFET L=6.4e-08
+ W=5.6e-07 AD=6.328e-14 AS=1.2768e-13 PD=7.86e-07 PS=1.016e-06 NRD=0.201786
+ NRS=0.408929 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=4.698e-06
+ SB=1.203e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.256e-15 PANW10=2.7584e-14
XMMN10 N_E_MMN10_d N_C_MMN10_g N_VSS_MMN12_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.6e-07 AD=1.2712e-13 AS=1.2768e-13 PD=1.014e-06 PS=1.016e-06
+ NRD=0.371429 NRS=0.405357 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=5e-06 SB=6.82e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN11 N_E_MMN10_d N_R_MMN11_g N_VSS_MMN11_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.6e-07 AD=1.2712e-13 AS=9.128e-14 PD=1.014e-06 PS=1.446e-06
+ NRD=0.439286 NRS=0.180357 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=5e-06 SB=1.63e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN14 N_Q_MMN14_d N_C_MMN14_g N_VSS_MMN14_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.6e-07 AD=1.4336e-13 AS=1.1144e-13 PD=1.632e-06 PS=1.518e-06
+ NRD=0.348214 NRS=0.180357 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.99e-07 SB=2.56e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMP0 N_CLK-_MMP0_d N_CLK_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.55e-07 AD=1.6426e-13 AS=2.14397e-13 PD=2.254e-06 PS=1.404e-06
+ NRD=0.108901 NRS=0.363351 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.72e-07 SB=6.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=4.011e-14
+ PANW6=2.1965e-14 PANW7=0 PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP1 N_CLK+_MMP1_d N_CLK-_MMP1_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.55e-07 AD=1.61395e-13 AS=2.14397e-13 PD=2.248e-06 PS=1.404e-06
+ NRD=0.105759 NRS=0.106806 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=6.86e-07 SB=1.69e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=2.947e-14 PANW9=6.4195e-14 PANW10=7.2345e-14
XMMP4 N_B_MMP4_d N_R_MMP4_g NET6 N_VDD_D0_noxref_neg PFET L=6.5e-08 W=9.55e-07
+ AD=1.5853e-13 AS=2.37795e-13 PD=2.242e-06 PS=1.453e-06 NRD=0.10555
+ NRS=0.260733 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.66e-07
+ SB=5e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=2.886e-14 PANW10=1.3442e-13
XMMP5 NET6 N_A_MMP5_g N_VDD_MMP5_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.37795e-13 AS=2.17262e-13 PD=1.453e-06 PS=1.41e-06 NRD=0.260733
+ NRS=0.232461 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=7.29e-07
+ SB=5e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP2 NET5 N_D_MMP2_g N_VDD_MMP5_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.32542e-13 AS=2.17262e-13 PD=1.442e-06 PS=1.41e-06 NRD=0.254974
+ NRS=0.243979 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.249e-06
+ SB=4.651e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP3 N_A_MMP3_d N_CLK+_MMP3_g NET5 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.18217e-13 AS=2.32542e-13 PD=1.412e-06 PS=1.442e-06
+ NRD=0.208377 NRS=0.254974 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.801e-06 SB=4.099e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP7 N_A_MMP3_d N_CLK-_MMP7_g NET7 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.18217e-13 AS=2.18695e-13 PD=1.412e-06 PS=1.413e-06
+ NRD=0.270157 NRS=0.239791 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=2.323e-06 SB=3.577e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP6 NET7 N_B_MMP6_g N_VDD_MMP6_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.18695e-13 AS=2.17262e-13 PD=1.413e-06 PS=1.41e-06 NRD=0.239791
+ NRS=0.248168 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.846e-06
+ SB=3.054e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP8 NET8 N_B_MMP8_g N_VDD_MMP6_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.17262e-13 AS=2.17262e-13 PD=1.41e-06 PS=1.41e-06 NRD=0.23822
+ NRS=0.228272 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.366e-06
+ SB=2.534e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP9 N_C_MMP9_d N_CLK-_MMP9_g NET8 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.1774e-13 AS=2.17262e-13 PD=1.411e-06 PS=1.41e-06 NRD=0.224084
+ NRS=0.23822 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.886e-06
+ SB=2.014e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP13 N_C_MMP9_d N_CLK+_MMP13_g NET10 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.1774e-13 AS=1.07915e-13 PD=1.411e-06 PS=1.181e-06 NRD=0.253403
+ NRS=0.118325 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.407e-06
+ SB=1.493e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP12 NET10 N_E_MMP12_g N_VDD_MMP12_s N_VDD_D0_noxref_neg PFET L=6.4e-08
+ W=9.55e-07 AD=1.07915e-13 AS=2.1774e-13 PD=1.181e-06 PS=1.411e-06 NRD=0.118325
+ NRS=0.224084 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.698e-06
+ SB=1.203e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.688e-15 PANW9=2.8416e-14 PANW10=7.1232e-14
XMMP11 NET9 N_C_MMP11_g N_VDD_MMP12_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.16785e-13 AS=2.1774e-13 PD=1.409e-06 PS=1.411e-06 NRD=0.237696
+ NRS=0.253403 M=1 NF=1 CNR_SWITCH=2 PCCRIT=0 PAR=1 PTWELL=1 SA=5e-06
+ SB=6.82e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=2.886e-14 PANW10=1.3442e-13
XMMP10 N_E_MMP10_d N_R_MMP10_g NET9 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=1.55665e-13 AS=2.16785e-13 PD=2.236e-06 PS=1.409e-06
+ NRD=0.104712 NRS=0.237696 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=5e-06 SB=1.63e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=2.73e-15 PANW9=9.0935e-14 PANW10=7.2345e-14
XMMP14 N_Q_MMP14_d N_C_MMP14_g N_VDD_MMP14_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.55e-07 AD=2.4448e-13 AS=1.90045e-13 PD=2.422e-06 PS=2.308e-06
+ NRD=0.19267 NRS=0.114136 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.99e-07 SB=2.56e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=6.2075e-14 PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
*
.include "DFF.pex.sp.DFF.pxi"
*
.ends
*
*
