* File: nand2.pex.sp
* Created: Tue Apr 15 11:58:04 2025
* Program "Calibre xRC"
* Version "v2024.4_12.9"
*
.include "nand2.pex.sp.pex"
.subckt nand2  OUT GND! VDD! INA INB
* 
* INB	INB
* INA	INA
* VDD!	VDD!
* GND!	GND!
* OUT	OUT
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=5.67424e-12
+ PERIM=9.616e-06
XMMN0 N_OUT_MMN0_d N_INA_MMN0_g NET1 N_GND!_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=9.296e-14 AS=2.1644e-13 PD=1.452e-06 PS=1.333e-06 NRD=0.183929
+ NRS=0.690179 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.66e-07
+ SB=1.267e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=1.1505e-14 PANW9=2.4895e-14 PANW10=0
XMMN1 NET1 N_INB_MMN1_g N_GND!_MMN1_s N_GND!_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=2.1644e-13 AS=2.4024e-13 PD=1.333e-06 PS=1.978e-06 NRD=0.690179
+ NRS=0.624405 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.004e-06
+ SB=4.29e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=1.1505e-14 PANW9=2.4895e-14 PANW10=0
XMMP0 N_OUT_MMP0_d N_INA_MMP0_g N_VDD!_MMP0_s N_VDD!_D0_noxref_neg PFET
+ L=6.5e-08 W=9.55e-07 AD=1.5853e-13 AS=3.69107e-13 PD=2.242e-06 PS=1.728e-06
+ NRD=0.110995 NRS=0.238743 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.66e-07 SB=1.267e-06 SD=0 PANW1=4.615e-15 PANW2=3.25e-15 PANW3=3.25e-15
+ PANW4=4.205e-15 PANW5=5.1e-14 PANW6=1.987e-14 PANW7=1.3e-14 PANW8=1.3e-14
+ PANW9=1.196e-14 PANW10=9.1715e-14
XMMP1 N_OUT_MMP1_d N_INB_MMP1_g N_VDD!_MMP0_s N_VDD!_D0_noxref_neg PFET
+ L=6.5e-08 W=9.55e-07 AD=4.09695e-13 AS=3.69107e-13 PD=2.768e-06 PS=1.728e-06
+ NRD=0.376963 NRS=0.570681 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.004e-06 SB=4.29e-07 SD=0 PANW1=4.615e-15 PANW2=3.25e-15 PANW3=3.25e-15
+ PANW4=3.25e-15 PANW5=3.25e-15 PANW6=6.5e-15 PANW7=7.5075e-14 PANW8=1.3e-14
+ PANW9=7.4035e-14 PANW10=2.964e-14
*
.include "nand2.pex.sp.NAND2.pxi"
*
.ends
*
*
