* File: XNOR2.pex.sp
* Created: Thu May  8 20:46:51 2025
* Program "Calibre xRC"
* Version "v2024.4_12.9"
* 
.include "XNOR2.pex.sp.pex"
.subckt XNOR2  VSS OUT VDD A B
* 
* B	B
* A	A
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=9.34934e-12
+ PERIM=1.2258e-05
XMMN0 N_Z_MMN0_d N_A_MMN0_g NET1 N_VSS_D0_noxref_pos NFET L=6.5e-08 W=5.6e-07
+ AD=9.296e-14 AS=1.386e-13 PD=1.452e-06 PS=1.055e-06 NRD=0.178571 NRS=0.441964
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.66e-07 SB=2.038e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0
+ PANW9=8.385e-15 PANW10=2.8015e-14
XMMN1 NET1 N_B_MMN1_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.386e-13 AS=9.772e-14 PD=1.055e-06 PS=9.09e-07 NRD=0.441964
+ NRS=0.178571 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=7.26e-07
+ SB=1.478e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN4 N_NET3_MMN4_d N_Z_MMN4_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=9.1e-14 AS=9.772e-14 PD=8.85e-07 PS=9.09e-07 NRD=0.394643
+ NRS=0.444643 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.14e-06
+ SB=1.064e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN3 N_OUT_MMN3_d N_B_MMN3_g N_NET3_MMN4_d N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.232e-13 AS=9.1e-14 PD=1e-06 PS=8.85e-07 NRD=0.605357
+ NRS=0.185714 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.53e-06
+ SB=6.74e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMN2 N_OUT_MMN3_d N_A_MMN2_g N_NET3_MMN2_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.232e-13 AS=9.464e-14 PD=1e-06 PS=1.458e-06 NRD=0.180357
+ NRS=0.183929 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.035e-06
+ SB=1.69e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=8.385e-15 PANW10=2.8015e-14
XMMP0 N_Z_MMP0_d N_A_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.36362e-13 AS=1.5853e-13 PD=1.45e-06 PS=2.242e-06 NRD=0.127749
+ NRS=0.106806 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.66e-07
+ SB=2.038e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=1.6235e-14 PANW5=4.584e-14
+ PANW6=0 PANW7=0 PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
XMMP1 N_Z_MMP0_d N_B_MMP1_g N_VDD_MMP1_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.36362e-13 AS=1.66647e-13 PD=1.45e-06 PS=1.304e-06 NRD=0.390576
+ NRS=0.12356 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=7.26e-07
+ SB=1.478e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=9.415e-15 PANW9=8.425e-14 PANW10=1.3442e-13
XMMP4 N_OUT_MMP4_d N_Z_MMP4_g N_VDD_MMP1_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=1.55187e-13 AS=1.66647e-13 PD=1.28e-06 PS=1.304e-06 NRD=0.230366
+ NRS=0.241885 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.14e-06
+ SB=1.064e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=2.73e-15 PANW9=4.032e-14 PANW10=1.85035e-13
XMMP2 N_OUT_MMP4_d N_B_MMP2_g NET2 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=1.55187e-13 AS=2.101e-13 PD=1.28e-06 PS=1.395e-06 NRD=0.109948
+ NRS=0.230366 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.53e-06
+ SB=6.74e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=4.64e-15 PANW9=8.9025e-14 PANW10=1.3442e-13
XMMP3 NET2 N_A_MMP3_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.55e-07 AD=2.101e-13 AS=1.61395e-13 PD=1.395e-06 PS=2.248e-06 NRD=0.230366
+ NRS=0.104712 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.035e-06
+ SB=1.69e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=6.685e-15
+ PANW6=5.539e-14 PANW7=0 PANW8=2.73e-15 PANW9=2.886e-14 PANW10=7.2345e-14
*
.include "XNOR2.pex.sp.XNOR2.pxi"
*
.ends
*
*
