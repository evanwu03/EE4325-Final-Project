// Created by ihdl
module UART (
	i_System_Clock, 
	i_Rst_L, 
	i_TX_Valid, 
	i_TX_Byte, 
	i_RX_Serial, 
	o_TX_Busy, 
	o_TX_Serial, 
	o_TX_Done, 
	o_RX_Done, 
	o_RX_Byte);
   input i_System_Clock;
   input i_Rst_L;
   input i_TX_Valid;
   input [7:0] i_TX_Byte;
   input i_RX_Serial;
   output o_TX_Busy;
   output o_TX_Serial;
   output o_TX_Done;
   output o_RX_Done;
   output [7:0] o_RX_Byte;

   // Internal wires
   wire \UART_RX_Inst/n168 ;
   wire \UART_RX_Inst/n167 ;
   wire \UART_RX_Inst/n166 ;
   wire \UART_RX_Inst/n165 ;
   wire \UART_RX_Inst/n164 ;
   wire \UART_RX_Inst/n163 ;
   wire \UART_RX_Inst/n162 ;
   wire \UART_RX_Inst/n161 ;
   wire \UART_RX_Inst/n160 ;
   wire \UART_RX_Inst/n159 ;
   wire \UART_RX_Inst/n158 ;
   wire \UART_RX_Inst/n157 ;
   wire \UART_RX_Inst/n156 ;
   wire \UART_RX_Inst/n155 ;
   wire \UART_RX_Inst/n154 ;
   wire \UART_RX_Inst/n153 ;
   wire \UART_RX_Inst/n152 ;
   wire \UART_RX_Inst/n151 ;
   wire \UART_RX_Inst/n150 ;
   wire \UART_RX_Inst/n149 ;
   wire \UART_RX_Inst/n148 ;
   wire \UART_RX_Inst/n147 ;
   wire \UART_RX_Inst/n146 ;
   wire \UART_RX_Inst/n145 ;
   wire \UART_RX_Inst/n144 ;
   wire \UART_RX_Inst/n143 ;
   wire \UART_RX_Inst/n142 ;
   wire \UART_RX_Inst/n141 ;
   wire \UART_RX_Inst/n140 ;
   wire \UART_RX_Inst/n139 ;
   wire \UART_RX_Inst/n138 ;
   wire \UART_RX_Inst/n137 ;
   wire \UART_RX_Inst/n136 ;
   wire \UART_RX_Inst/n135 ;
   wire \UART_RX_Inst/n134 ;
   wire \UART_RX_Inst/n133 ;
   wire \UART_RX_Inst/n132 ;
   wire \UART_RX_Inst/n131 ;
   wire \UART_RX_Inst/n130 ;
   wire \UART_RX_Inst/n129 ;
   wire \UART_RX_Inst/n128 ;
   wire \UART_RX_Inst/n127 ;
   wire \UART_RX_Inst/n126 ;
   wire \UART_RX_Inst/n125 ;
   wire \UART_RX_Inst/n124 ;
   wire \UART_RX_Inst/n123 ;
   wire \UART_RX_Inst/n122 ;
   wire \UART_RX_Inst/n121 ;
   wire \UART_RX_Inst/n120 ;
   wire \UART_RX_Inst/n119 ;
   wire \UART_RX_Inst/n118 ;
   wire \UART_RX_Inst/n117 ;
   wire \UART_RX_Inst/n116 ;
   wire \UART_RX_Inst/n115 ;
   wire \UART_RX_Inst/n114 ;
   wire \UART_RX_Inst/n113 ;
   wire \UART_RX_Inst/n112 ;
   wire \UART_RX_Inst/n111 ;
   wire \UART_RX_Inst/n110 ;
   wire \UART_RX_Inst/n109 ;
   wire \UART_RX_Inst/n108 ;
   wire \UART_RX_Inst/n107 ;
   wire \UART_RX_Inst/n106 ;
   wire \UART_RX_Inst/n105 ;
   wire \UART_RX_Inst/n104 ;
   wire \UART_RX_Inst/n103 ;
   wire \UART_RX_Inst/n102 ;
   wire \UART_RX_Inst/n101 ;
   wire \UART_RX_Inst/n100 ;
   wire \UART_RX_Inst/n99 ;
   wire \UART_RX_Inst/n98 ;
   wire \UART_RX_Inst/n97 ;
   wire \UART_RX_Inst/n96 ;
   wire \UART_RX_Inst/n95 ;
   wire \UART_RX_Inst/n94 ;
   wire \UART_RX_Inst/n93 ;
   wire \UART_RX_Inst/n92 ;
   wire \UART_RX_Inst/n91 ;
   wire \UART_RX_Inst/n90 ;
   wire \UART_RX_Inst/n89 ;
   wire \UART_RX_Inst/n88 ;
   wire \UART_RX_Inst/n87 ;
   wire \UART_RX_Inst/n86 ;
   wire \UART_RX_Inst/n85 ;
   wire \UART_RX_Inst/n84 ;
   wire \UART_RX_Inst/n83 ;
   wire \UART_RX_Inst/n82 ;
   wire \UART_RX_Inst/n81 ;
   wire \UART_RX_Inst/n80 ;
   wire \UART_RX_Inst/n79 ;
   wire \UART_RX_Inst/n78 ;
   wire \UART_RX_Inst/n77 ;
   wire \UART_RX_Inst/n76 ;
   wire \UART_RX_Inst/n75 ;
   wire \UART_RX_Inst/n73 ;
   wire \UART_RX_Inst/n72 ;
   wire \UART_RX_Inst/n71 ;
   wire \UART_RX_Inst/n70 ;
   wire \UART_RX_Inst/n69 ;
   wire \UART_RX_Inst/n68 ;
   wire \UART_RX_Inst/n67 ;
   wire \UART_RX_Inst/n66 ;
   wire \UART_RX_Inst/n65 ;
   wire \UART_RX_Inst/n64 ;
   wire \UART_RX_Inst/n63 ;
   wire \UART_RX_Inst/n62 ;
   wire \UART_RX_Inst/n61 ;
   wire \UART_RX_Inst/n60 ;
   wire \UART_RX_Inst/n59 ;
   wire \UART_RX_Inst/n58 ;
   wire \UART_RX_Inst/n57 ;
   wire \UART_RX_Inst/n56 ;
   wire \UART_RX_Inst/n55 ;
   wire \UART_RX_Inst/n54 ;
   wire \UART_RX_Inst/n53 ;
   wire \UART_RX_Inst/n52 ;
   wire \UART_RX_Inst/n51 ;
   wire \UART_RX_Inst/n50 ;
   wire \UART_RX_Inst/n49 ;
   wire \UART_RX_Inst/n48 ;
   wire \UART_RX_Inst/n47 ;
   wire \UART_RX_Inst/n46 ;
   wire \UART_RX_Inst/n45 ;
   wire \UART_RX_Inst/n44 ;
   wire \UART_RX_Inst/n43 ;
   wire \UART_RX_Inst/n42 ;
   wire \UART_RX_Inst/n41 ;
   wire \UART_RX_Inst/n40 ;
   wire \UART_RX_Inst/n39 ;
   wire \UART_RX_Inst/n38 ;
   wire \UART_RX_Inst/n37 ;
   wire \UART_RX_Inst/n36 ;
   wire \UART_RX_Inst/n35 ;
   wire \UART_RX_Inst/n34 ;
   wire \UART_RX_Inst/n33 ;
   wire \UART_RX_Inst/n32 ;
   wire \UART_RX_Inst/n31 ;
   wire \UART_RX_Inst/n30 ;
   wire \UART_RX_Inst/n29 ;
   wire \UART_RX_Inst/n28 ;
   wire \UART_RX_Inst/n27 ;
   wire \UART_RX_Inst/n26 ;
   wire \UART_RX_Inst/n25 ;
   wire \UART_RX_Inst/n24 ;
   wire \UART_RX_Inst/n23 ;
   wire \UART_RX_Inst/n22 ;
   wire \UART_RX_Inst/n21 ;
   wire \UART_RX_Inst/n20 ;
   wire \UART_RX_Inst/n19 ;
   wire \UART_RX_Inst/n18 ;
   wire \UART_RX_Inst/n17 ;
   wire \UART_RX_Inst/n16 ;
   wire \UART_RX_Inst/U3/U1/Z_9 ;
   wire \UART_RX_Inst/U3/U1/Z_7 ;
   wire \UART_RX_Inst/N226 ;
   wire \UART_RX_Inst/N225 ;
   wire \UART_RX_Inst/N224 ;
   wire \UART_RX_Inst/N223 ;
   wire \UART_RX_Inst/N222 ;
   wire \UART_RX_Inst/N221 ;
   wire \UART_RX_Inst/N220 ;
   wire \UART_RX_Inst/N219 ;
   wire \UART_RX_Inst/N213 ;
   wire \UART_RX_Inst/N212 ;
   wire \UART_RX_Inst/N211 ;
   wire \UART_RX_Inst/N210 ;
   wire \UART_RX_Inst/N209 ;
   wire \UART_RX_Inst/N208 ;
   wire \UART_RX_Inst/N207 ;
   wire \UART_RX_Inst/N206 ;
   wire \UART_RX_Inst/N205 ;
   wire \UART_RX_Inst/N204 ;
   wire \UART_RX_Inst/N203 ;
   wire \UART_RX_Inst/N202 ;
   wire \UART_RX_Inst/N201 ;
   wire \UART_RX_Inst/N200 ;
   wire \UART_RX_Inst/N199 ;
   wire \UART_RX_Inst/N198 ;
   wire \UART_RX_Inst/N197 ;
   wire \UART_RX_Inst/N196 ;
   wire \UART_RX_Inst/N195 ;
   wire \UART_RX_Inst/N194 ;
   wire \UART_RX_Inst/N193 ;
   wire \UART_RX_Inst/N192 ;
   wire \UART_RX_Inst/N191 ;
   wire \UART_RX_Inst/N190 ;
   wire \UART_RX_Inst/N189 ;
   wire \UART_RX_Inst/N188 ;
   wire \UART_RX_Inst/N187 ;
   wire \UART_RX_Inst/N186 ;
   wire \UART_RX_Inst/N185 ;
   wire \UART_RX_Inst/N184 ;
   wire \UART_RX_Inst/N183 ;
   wire \UART_RX_Inst/N182 ;
   wire \UART_RX_Inst/N181 ;
   wire \UART_RX_Inst/N180 ;
   wire \UART_RX_Inst/N145 ;
   wire \UART_RX_Inst/N114 ;
   wire \UART_RX_Inst/N113 ;
   wire \UART_RX_Inst/N112 ;
   wire \UART_RX_Inst/N102 ;
   wire \UART_RX_Inst/N101 ;
   wire \UART_RX_Inst/N100 ;
   wire \UART_RX_Inst/N99 ;
   wire \UART_RX_Inst/N98 ;
   wire \UART_RX_Inst/N97 ;
   wire \UART_RX_Inst/N96 ;
   wire \UART_RX_Inst/N95 ;
   wire \UART_RX_Inst/N94 ;
   wire \UART_RX_Inst/N93 ;
   wire \UART_RX_Inst/N92 ;
   wire \UART_RX_Inst/N91 ;
   wire \UART_RX_Inst/N90 ;
   wire \UART_RX_Inst/N89 ;
   wire \UART_RX_Inst/N88 ;
   wire \UART_RX_Inst/N87 ;
   wire \UART_RX_Inst/N84 ;
   wire \UART_RX_Inst/N39 ;
   wire \UART_RX_Inst/N38 ;
   wire \UART_RX_Inst/N37 ;
   wire \UART_RX_Inst/N35 ;
   wire \UART_RX_Inst/N34 ;
   wire \UART_RX_Inst/N33 ;
   wire \UART_RX_Inst/N32 ;
   wire \UART_RX_Inst/N31 ;
   wire \UART_RX_Inst/N29 ;
   wire \UART_RX_Inst/N28 ;
   wire \UART_RX_Inst/N26 ;
   wire \UART_RX_Inst/N24 ;
   wire \UART_RX_Inst/N23 ;
   wire \UART_RX_Inst/N21 ;
   wire \UART_RX_Inst/r_Bit_Index[0] ;
   wire \UART_RX_Inst/N11 ;
   wire \UART_RX_Inst/N10 ;
   wire \UART_RX_Inst/N9 ;
   wire \UART_RX_Inst/N8 ;
   wire \UART_RX_Inst/N7 ;
   wire \UART_RX_Inst/N6 ;
   wire \UART_RX_Inst/N5 ;
   wire \UART_RX_Inst/N4 ;
   wire \UART_RX_Inst/N3 ;
   wire \UART_RX_Inst/N2 ;
   wire \UART_RX_Inst/N1 ;
   wire \UART_RX_Inst/N0 ;
   wire \UART_TX_Inst/n122 ;
   wire \UART_TX_Inst/n121 ;
   wire \UART_TX_Inst/n120 ;
   wire \UART_TX_Inst/n119 ;
   wire \UART_TX_Inst/n118 ;
   wire \UART_TX_Inst/n117 ;
   wire \UART_TX_Inst/n116 ;
   wire \UART_TX_Inst/n115 ;
   wire \UART_TX_Inst/n114 ;
   wire \UART_TX_Inst/n113 ;
   wire \UART_TX_Inst/n112 ;
   wire \UART_TX_Inst/n111 ;
   wire \UART_TX_Inst/n110 ;
   wire \UART_TX_Inst/n109 ;
   wire \UART_TX_Inst/n108 ;
   wire \UART_TX_Inst/n107 ;
   wire \UART_TX_Inst/n106 ;
   wire \UART_TX_Inst/n105 ;
   wire \UART_TX_Inst/n104 ;
   wire \UART_TX_Inst/n103 ;
   wire \UART_TX_Inst/n102 ;
   wire \UART_TX_Inst/n101 ;
   wire \UART_TX_Inst/n100 ;
   wire \UART_TX_Inst/n99 ;
   wire \UART_TX_Inst/n98 ;
   wire \UART_TX_Inst/n97 ;
   wire \UART_TX_Inst/n96 ;
   wire \UART_TX_Inst/n95 ;
   wire \UART_TX_Inst/n94 ;
   wire \UART_TX_Inst/n93 ;
   wire \UART_TX_Inst/n92 ;
   wire \UART_TX_Inst/n91 ;
   wire \UART_TX_Inst/n90 ;
   wire \UART_TX_Inst/n89 ;
   wire \UART_TX_Inst/n88 ;
   wire \UART_TX_Inst/n87 ;
   wire \UART_TX_Inst/n86 ;
   wire \UART_TX_Inst/n85 ;
   wire \UART_TX_Inst/n84 ;
   wire \UART_TX_Inst/n83 ;
   wire \UART_TX_Inst/n82 ;
   wire \UART_TX_Inst/n81 ;
   wire \UART_TX_Inst/n80 ;
   wire \UART_TX_Inst/n79 ;
   wire \UART_TX_Inst/n78 ;
   wire \UART_TX_Inst/n77 ;
   wire \UART_TX_Inst/n76 ;
   wire \UART_TX_Inst/n75 ;
   wire \UART_TX_Inst/n74 ;
   wire \UART_TX_Inst/n73 ;
   wire \UART_TX_Inst/n72 ;
   wire \UART_TX_Inst/n71 ;
   wire \UART_TX_Inst/n70 ;
   wire \UART_TX_Inst/n69 ;
   wire \UART_TX_Inst/n68 ;
   wire \UART_TX_Inst/n67 ;
   wire \UART_TX_Inst/n66 ;
   wire \UART_TX_Inst/n65 ;
   wire \UART_TX_Inst/n64 ;
   wire \UART_TX_Inst/n63 ;
   wire \UART_TX_Inst/n62 ;
   wire \UART_TX_Inst/n61 ;
   wire \UART_TX_Inst/n60 ;
   wire \UART_TX_Inst/n59 ;
   wire \UART_TX_Inst/n58 ;
   wire \UART_TX_Inst/n57 ;
   wire \UART_TX_Inst/n56 ;
   wire \UART_TX_Inst/n55 ;
   wire \UART_TX_Inst/n54 ;
   wire \UART_TX_Inst/n53 ;
   wire \UART_TX_Inst/n52 ;
   wire \UART_TX_Inst/n51 ;
   wire \UART_TX_Inst/n50 ;
   wire \UART_TX_Inst/n49 ;
   wire \UART_TX_Inst/n48 ;
   wire \UART_TX_Inst/n47 ;
   wire \UART_TX_Inst/n46 ;
   wire \UART_TX_Inst/n45 ;
   wire \UART_TX_Inst/n44 ;
   wire \UART_TX_Inst/n43 ;
   wire \UART_TX_Inst/n42 ;
   wire \UART_TX_Inst/n41 ;
   wire \UART_TX_Inst/n39 ;
   wire \UART_TX_Inst/n37 ;
   wire \UART_TX_Inst/n36 ;
   wire \UART_TX_Inst/n35 ;
   wire \UART_TX_Inst/n34 ;
   wire \UART_TX_Inst/n33 ;
   wire \UART_TX_Inst/n32 ;
   wire \UART_TX_Inst/n31 ;
   wire \UART_TX_Inst/n30 ;
   wire \UART_TX_Inst/n29 ;
   wire \UART_TX_Inst/n28 ;
   wire \UART_TX_Inst/n27 ;
   wire \UART_TX_Inst/n26 ;
   wire \UART_TX_Inst/n25 ;
   wire \UART_TX_Inst/n24 ;
   wire \UART_TX_Inst/n23 ;
   wire \UART_TX_Inst/n22 ;
   wire \UART_TX_Inst/n21 ;
   wire \UART_TX_Inst/n20 ;
   wire \UART_TX_Inst/n19 ;
   wire \UART_TX_Inst/n18 ;
   wire \UART_TX_Inst/n17 ;
   wire \UART_TX_Inst/n16 ;
   wire \UART_TX_Inst/n15 ;
   wire \UART_TX_Inst/n14 ;
   wire \UART_TX_Inst/n13 ;
   wire \UART_TX_Inst/n12 ;
   wire \UART_TX_Inst/n11 ;
   wire \UART_TX_Inst/n10 ;
   wire \UART_TX_Inst/n9 ;
   wire \UART_TX_Inst/n8 ;
   wire \UART_TX_Inst/N146 ;
   wire \UART_TX_Inst/N145 ;
   wire \UART_TX_Inst/N144 ;
   wire \UART_TX_Inst/N143 ;
   wire \UART_TX_Inst/N142 ;
   wire \UART_TX_Inst/N141 ;
   wire \UART_TX_Inst/N140 ;
   wire \UART_TX_Inst/N139 ;
   wire \UART_TX_Inst/N138 ;
   wire \UART_TX_Inst/N137 ;
   wire \UART_TX_Inst/N136 ;
   wire \UART_TX_Inst/N129 ;
   wire \UART_TX_Inst/N127 ;
   wire \UART_TX_Inst/N126 ;
   wire \UART_TX_Inst/N125 ;
   wire \UART_TX_Inst/N124 ;
   wire \UART_TX_Inst/N123 ;
   wire \UART_TX_Inst/N122 ;
   wire \UART_TX_Inst/N121 ;
   wire \UART_TX_Inst/N120 ;
   wire \UART_TX_Inst/N119 ;
   wire \UART_TX_Inst/N118 ;
   wire \UART_TX_Inst/N117 ;
   wire \UART_TX_Inst/N116 ;
   wire \UART_TX_Inst/N115 ;
   wire \UART_TX_Inst/N114 ;
   wire \UART_TX_Inst/N113 ;
   wire \UART_TX_Inst/N112 ;
   wire \UART_TX_Inst/N111 ;
   wire \UART_TX_Inst/N110 ;
   wire \UART_TX_Inst/N97 ;
   wire \UART_TX_Inst/N96 ;
   wire \UART_TX_Inst/N95 ;
   wire \UART_TX_Inst/N94 ;
   wire \UART_TX_Inst/N93 ;
   wire \UART_TX_Inst/N92 ;
   wire \UART_TX_Inst/N91 ;
   wire \UART_TX_Inst/N90 ;
   wire \UART_TX_Inst/N89 ;
   wire \UART_TX_Inst/N88 ;
   wire \UART_TX_Inst/N87 ;
   wire \UART_TX_Inst/N68 ;
   wire \UART_TX_Inst/N67 ;
   wire \UART_TX_Inst/N66 ;
   wire \UART_TX_Inst/N64 ;
   wire \UART_TX_Inst/N23 ;
   wire \UART_TX_Inst/N20 ;
   wire \UART_TX_Inst/N18 ;
   wire \UART_TX_Inst/N17 ;
   wire \UART_TX_Inst/N16 ;
   wire \UART_TX_Inst/N12 ;
   wire \UART_TX_Inst/N9 ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire [2:1] \UART_RX_Inst/lt_110/LTV ;
   wire [2:0] \UART_RX_Inst/lt_110/AEQB ;
   wire [2:0] \UART_RX_Inst/lt_110/LTV1 ;
   wire [2:0] \UART_RX_Inst/lt_110/LTV2 ;
   wire [15:0] \UART_RX_Inst/r_Clock_Count ;
   wire [2:0] \UART_RX_Inst/r_RX_State ;
   wire [2:1] \UART_TX_Inst/lt_109/LTV ;
   wire [2:0] \UART_TX_Inst/lt_109/AEQB ;
   wire [2:0] \UART_TX_Inst/lt_109/LTV1 ;
   wire [2:0] \UART_TX_Inst/lt_109/LTV2 ;
   wire [7:0] \UART_TX_Inst/r_TX_Data ;
   wire [10:0] \UART_TX_Inst/r_Clock_Count ;
   wire [1:0] \UART_TX_Inst/r_SM_Main ;
   wire [10:0] \UART_TX_Inst/r31/LTV2 ;
   wire [10:0] \UART_TX_Inst/r31/LTV1 ;
   wire [10:0] \UART_TX_Inst/r31/AEQB ;
   wire [10:1] \UART_TX_Inst/r31/LTV ;
   wire [15:0] \UART_RX_Inst/r35/LTV2 ;
   wire [15:0] \UART_RX_Inst/r35/LTV1 ;
   wire [15:0] \UART_RX_Inst/r35/AEQB ;
   wire [15:1] \UART_RX_Inst/r35/LTV ;

   INV \UART_RX_Inst/U193  (.OUT(\UART_RX_Inst/n168 ),
	.IN(\UART_RX_Inst/r_Bit_Index[0] ));
   INV \UART_RX_Inst/U192  (.OUT(\UART_RX_Inst/n167 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [1]));
   INV \UART_RX_Inst/U187  (.OUT(\UART_RX_Inst/N226 ),
	.IN(\UART_RX_Inst/n137 ));
   INV \UART_RX_Inst/U186  (.OUT(\UART_RX_Inst/N225 ),
	.IN(\UART_RX_Inst/n136 ));
   INV \UART_RX_Inst/U185  (.OUT(\UART_RX_Inst/N224 ),
	.IN(\UART_RX_Inst/n135 ));
   INV \UART_RX_Inst/U184  (.OUT(\UART_RX_Inst/N223 ),
	.IN(\UART_RX_Inst/n134 ));
   INV \UART_RX_Inst/U183  (.OUT(\UART_RX_Inst/N222 ),
	.IN(\UART_RX_Inst/n133 ));
   INV \UART_RX_Inst/U182  (.OUT(\UART_RX_Inst/N221 ),
	.IN(\UART_RX_Inst/n132 ));
   INV \UART_RX_Inst/U181  (.OUT(\UART_RX_Inst/N220 ),
	.IN(\UART_RX_Inst/n131 ));
   INV \UART_RX_Inst/U180  (.OUT(\UART_RX_Inst/N219 ),
	.IN(\UART_RX_Inst/n130 ));
   INV \UART_RX_Inst/U179  (.OUT(\UART_RX_Inst/N26 ),
	.IN(\UART_RX_Inst/n83 ));
   INV \UART_RX_Inst/U178  (.OUT(\UART_RX_Inst/n94 ),
	.IN(\UART_RX_Inst/N145 ));
   INV \UART_RX_Inst/U177  (.OUT(\UART_RX_Inst/n129 ),
	.IN(\UART_RX_Inst/N84 ));
   NAND3 \UART_RX_Inst/U176  (.OUT(\UART_RX_Inst/n97 ),
	.C(\UART_RX_Inst/N33 ),
	.B(\UART_RX_Inst/n129 ),
	.A(\UART_RX_Inst/n94 ));
   NAND3 \UART_RX_Inst/U175  (.OUT(\UART_RX_Inst/n89 ),
	.C(\UART_RX_Inst/N84 ),
	.B(\UART_RX_Inst/n94 ),
	.A(\UART_RX_Inst/N33 ));
   INV \UART_RX_Inst/U174  (.OUT(\UART_RX_Inst/n84 ),
	.IN(\UART_RX_Inst/r_RX_State [0]));
   NAND2 \UART_RX_Inst/U173  (.OUT(\UART_RX_Inst/n100 ),
	.B(\UART_RX_Inst/n84 ),
	.A(\UART_RX_Inst/N26 ));
   NAND3 \UART_RX_Inst/U172  (.OUT(\UART_RX_Inst/N180 ),
	.C(\UART_RX_Inst/n100 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n97 ));
   INV \UART_RX_Inst/U171  (.OUT(\UART_RX_Inst/n128 ),
	.IN(\UART_RX_Inst/N112 ));
   NOR2 \UART_RX_Inst/U170  (.OUT(\UART_RX_Inst/N181 ),
	.B(\UART_RX_Inst/n128 ),
	.A(\UART_RX_Inst/n89 ));
   INV \UART_RX_Inst/U169  (.OUT(\UART_RX_Inst/n127 ),
	.IN(\UART_RX_Inst/N113 ));
   NOR2 \UART_RX_Inst/U168  (.OUT(\UART_RX_Inst/N182 ),
	.B(\UART_RX_Inst/n127 ),
	.A(\UART_RX_Inst/n89 ));
   INV \UART_RX_Inst/U167  (.OUT(\UART_RX_Inst/n126 ),
	.IN(\UART_RX_Inst/N114 ));
   NOR2 \UART_RX_Inst/U166  (.OUT(\UART_RX_Inst/N183 ),
	.B(\UART_RX_Inst/n126 ),
	.A(\UART_RX_Inst/n89 ));
   INV \UART_RX_Inst/U165  (.OUT(\UART_RX_Inst/n102 ),
	.IN(\UART_RX_Inst/N202 ));
   INV \UART_RX_Inst/U164  (.OUT(\UART_RX_Inst/n92 ),
	.IN(\UART_RX_Inst/N33 ));
   NAND2 \UART_RX_Inst/U163  (.OUT(\UART_RX_Inst/U3/U1/Z_9 ),
	.B(\UART_RX_Inst/n92 ),
	.A(\UART_RX_Inst/n102 ));
   INV \UART_RX_Inst/U162  (.OUT(\UART_RX_Inst/n123 ),
	.IN(\UART_RX_Inst/U3/U1/Z_9 ));
   NAND2 \UART_RX_Inst/U161  (.OUT(\UART_RX_Inst/n125 ),
	.B(\UART_RX_Inst/n94 ),
	.A(i_RX_Serial));
   NAND2 \UART_RX_Inst/U160  (.OUT(\UART_RX_Inst/n124 ),
	.B(\UART_RX_Inst/n125 ),
	.A(\UART_RX_Inst/U3/U1/Z_7 ));
   NAND3 \UART_RX_Inst/U159  (.OUT(\UART_RX_Inst/N184 ),
	.C(\UART_RX_Inst/n124 ),
	.B(\UART_RX_Inst/n123 ),
	.A(\UART_RX_Inst/n100 ));
   INV \UART_RX_Inst/U158  (.OUT(\UART_RX_Inst/n103 ),
	.IN(\UART_RX_Inst/U3/U1/Z_7 ));
   NAND2 \UART_RX_Inst/U157  (.OUT(\UART_RX_Inst/n122 ),
	.B(\UART_RX_Inst/n103 ),
	.A(\UART_RX_Inst/n123 ));
   NAND2 \UART_RX_Inst/U156  (.OUT(\UART_RX_Inst/n105 ),
	.B(\UART_RX_Inst/n122 ),
	.A(\UART_RX_Inst/N145 ));
   INV \UART_RX_Inst/U155  (.OUT(\UART_RX_Inst/n121 ),
	.IN(\UART_RX_Inst/N87 ));
   NOR2 \UART_RX_Inst/U154  (.OUT(\UART_RX_Inst/N185 ),
	.B(\UART_RX_Inst/n121 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U153  (.OUT(\UART_RX_Inst/n120 ),
	.IN(\UART_RX_Inst/N88 ));
   NOR2 \UART_RX_Inst/U152  (.OUT(\UART_RX_Inst/N186 ),
	.B(\UART_RX_Inst/n120 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U151  (.OUT(\UART_RX_Inst/n119 ),
	.IN(\UART_RX_Inst/N89 ));
   NOR2 \UART_RX_Inst/U150  (.OUT(\UART_RX_Inst/N187 ),
	.B(\UART_RX_Inst/n119 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U149  (.OUT(\UART_RX_Inst/n118 ),
	.IN(\UART_RX_Inst/N90 ));
   NOR2 \UART_RX_Inst/U148  (.OUT(\UART_RX_Inst/N188 ),
	.B(\UART_RX_Inst/n118 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U147  (.OUT(\UART_RX_Inst/n117 ),
	.IN(\UART_RX_Inst/N91 ));
   NOR2 \UART_RX_Inst/U146  (.OUT(\UART_RX_Inst/N189 ),
	.B(\UART_RX_Inst/n117 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U145  (.OUT(\UART_RX_Inst/n116 ),
	.IN(\UART_RX_Inst/N92 ));
   NOR2 \UART_RX_Inst/U144  (.OUT(\UART_RX_Inst/N190 ),
	.B(\UART_RX_Inst/n116 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U143  (.OUT(\UART_RX_Inst/n115 ),
	.IN(\UART_RX_Inst/N93 ));
   NOR2 \UART_RX_Inst/U142  (.OUT(\UART_RX_Inst/N191 ),
	.B(\UART_RX_Inst/n115 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U141  (.OUT(\UART_RX_Inst/n114 ),
	.IN(\UART_RX_Inst/N94 ));
   NOR2 \UART_RX_Inst/U140  (.OUT(\UART_RX_Inst/N192 ),
	.B(\UART_RX_Inst/n114 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U139  (.OUT(\UART_RX_Inst/n113 ),
	.IN(\UART_RX_Inst/N95 ));
   NOR2 \UART_RX_Inst/U138  (.OUT(\UART_RX_Inst/N193 ),
	.B(\UART_RX_Inst/n113 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U137  (.OUT(\UART_RX_Inst/n112 ),
	.IN(\UART_RX_Inst/N96 ));
   NOR2 \UART_RX_Inst/U136  (.OUT(\UART_RX_Inst/N194 ),
	.B(\UART_RX_Inst/n112 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U135  (.OUT(\UART_RX_Inst/n111 ),
	.IN(\UART_RX_Inst/N97 ));
   NOR2 \UART_RX_Inst/U134  (.OUT(\UART_RX_Inst/N195 ),
	.B(\UART_RX_Inst/n111 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U133  (.OUT(\UART_RX_Inst/n110 ),
	.IN(\UART_RX_Inst/N98 ));
   NOR2 \UART_RX_Inst/U132  (.OUT(\UART_RX_Inst/N196 ),
	.B(\UART_RX_Inst/n110 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U131  (.OUT(\UART_RX_Inst/n109 ),
	.IN(\UART_RX_Inst/N99 ));
   NOR2 \UART_RX_Inst/U130  (.OUT(\UART_RX_Inst/N197 ),
	.B(\UART_RX_Inst/n109 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U129  (.OUT(\UART_RX_Inst/n108 ),
	.IN(\UART_RX_Inst/N100 ));
   NOR2 \UART_RX_Inst/U128  (.OUT(\UART_RX_Inst/N198 ),
	.B(\UART_RX_Inst/n108 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U127  (.OUT(\UART_RX_Inst/n107 ),
	.IN(\UART_RX_Inst/N101 ));
   NOR2 \UART_RX_Inst/U126  (.OUT(\UART_RX_Inst/N199 ),
	.B(\UART_RX_Inst/n107 ),
	.A(\UART_RX_Inst/n105 ));
   INV \UART_RX_Inst/U125  (.OUT(\UART_RX_Inst/n106 ),
	.IN(\UART_RX_Inst/N102 ));
   NOR2 \UART_RX_Inst/U124  (.OUT(\UART_RX_Inst/N200 ),
	.B(\UART_RX_Inst/n106 ),
	.A(\UART_RX_Inst/n105 ));
   NAND2 \UART_RX_Inst/U123  (.OUT(\UART_RX_Inst/n90 ),
	.B(\UART_RX_Inst/n94 ),
	.A(\UART_RX_Inst/N202 ));
   INV \UART_RX_Inst/U122  (.OUT(\UART_RX_Inst/n104 ),
	.IN(\UART_RX_Inst/N39 ));
   NAND3 \UART_RX_Inst/U121  (.OUT(\UART_RX_Inst/N201 ),
	.C(\UART_RX_Inst/n100 ),
	.B(\UART_RX_Inst/n104 ),
	.A(\UART_RX_Inst/n90 ));
   NAND2 \UART_RX_Inst/U120  (.OUT(\UART_RX_Inst/n101 ),
	.B(\UART_RX_Inst/n103 ),
	.A(\UART_RX_Inst/n102 ));
   NAND2 \UART_RX_Inst/U119  (.OUT(\UART_RX_Inst/n96 ),
	.B(\UART_RX_Inst/n101 ),
	.A(\UART_RX_Inst/N145 ));
   INV \UART_RX_Inst/U118  (.OUT(\UART_RX_Inst/n99 ),
	.IN(\UART_RX_Inst/n100 ));
   INV \UART_RX_Inst/U117  (.OUT(\UART_RX_Inst/n95 ),
	.IN(i_RX_Serial));
   NAND2 \UART_RX_Inst/U116  (.OUT(\UART_RX_Inst/n98 ),
	.B(\UART_RX_Inst/n95 ),
	.A(\UART_RX_Inst/n99 ));
   NAND3 \UART_RX_Inst/U115  (.OUT(\UART_RX_Inst/N203 ),
	.C(\UART_RX_Inst/n98 ),
	.B(\UART_RX_Inst/n97 ),
	.A(\UART_RX_Inst/n96 ));
   NAND3 \UART_RX_Inst/U114  (.OUT(\UART_RX_Inst/n91 ),
	.C(\UART_RX_Inst/U3/U1/Z_7 ),
	.B(\UART_RX_Inst/n95 ),
	.A(\UART_RX_Inst/n94 ));
   NAND2 \UART_RX_Inst/U113  (.OUT(\UART_RX_Inst/n93 ),
	.B(\UART_RX_Inst/N202 ),
	.A(\UART_RX_Inst/N145 ));
   NAND3 \UART_RX_Inst/U112  (.OUT(\UART_RX_Inst/N204 ),
	.C(\UART_RX_Inst/n93 ),
	.B(\UART_RX_Inst/n92 ),
	.A(\UART_RX_Inst/n91 ));
   INV \UART_RX_Inst/U111  (.OUT(\UART_RX_Inst/N205 ),
	.IN(\UART_RX_Inst/n90 ));
   NOR2 \UART_RX_Inst/U110  (.OUT(\UART_RX_Inst/N206 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n75 ));
   NOR2 \UART_RX_Inst/U109  (.OUT(\UART_RX_Inst/N207 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n76 ));
   NOR2 \UART_RX_Inst/U108  (.OUT(\UART_RX_Inst/N208 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n77 ));
   NOR2 \UART_RX_Inst/U107  (.OUT(\UART_RX_Inst/N209 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n78 ));
   NOR2 \UART_RX_Inst/U106  (.OUT(\UART_RX_Inst/N210 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n79 ));
   NOR2 \UART_RX_Inst/U105  (.OUT(\UART_RX_Inst/N211 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n80 ));
   NOR2 \UART_RX_Inst/U104  (.OUT(\UART_RX_Inst/N212 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n81 ));
   NOR2 \UART_RX_Inst/U103  (.OUT(\UART_RX_Inst/N213 ),
	.B(\UART_RX_Inst/n89 ),
	.A(\UART_RX_Inst/n82 ));
   INV \UART_RX_Inst/U102  (.OUT(\UART_RX_Inst/n88 ),
	.IN(\UART_RX_Inst/N28 ));
   NAND2 \UART_RX_Inst/U101  (.OUT(\UART_RX_Inst/N29 ),
	.B(\UART_RX_Inst/n88 ),
	.A(\UART_RX_Inst/r_RX_State [0]));
   NOR2 \UART_RX_Inst/U100  (.OUT(\UART_RX_Inst/n87 ),
	.B(\UART_RX_Inst/r_RX_State [0]),
	.A(\UART_RX_Inst/N31 ));
   INV \UART_RX_Inst/U99  (.OUT(\UART_RX_Inst/N32 ),
	.IN(\UART_RX_Inst/n87 ));
   INV \UART_RX_Inst/U98  (.OUT(\UART_RX_Inst/n86 ),
	.IN(\UART_RX_Inst/N34 ));
   NAND2 \UART_RX_Inst/U97  (.OUT(\UART_RX_Inst/N35 ),
	.B(\UART_RX_Inst/n86 ),
	.A(\UART_RX_Inst/r_RX_State [0]));
   NOR2 \UART_RX_Inst/U96  (.OUT(\UART_RX_Inst/n85 ),
	.B(\UART_RX_Inst/r_RX_State [0]),
	.A(\UART_RX_Inst/N37 ));
   INV \UART_RX_Inst/U95  (.OUT(\UART_RX_Inst/N38 ),
	.IN(\UART_RX_Inst/n85 ));
   INV \UART_RX_Inst/U93  (.OUT(\UART_RX_Inst/N112 ),
	.IN(\UART_RX_Inst/r_Bit_Index[0] ));
   INV \UART_RX_Inst/U92  (.OUT(\UART_RX_Inst/n65 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [1]));
   XNOR2 \UART_RX_Inst/U91  (.OUT(\UART_RX_Inst/N113 ),
	.B(\UART_RX_Inst/r_Bit_Index[0] ),
	.A(\UART_RX_Inst/n65 ));
   NAND2 \UART_RX_Inst/U90  (.OUT(\UART_RX_Inst/n73 ),
	.B(\UART_RX_Inst/r_Bit_Index[0] ),
	.A(\UART_RX_Inst/lt_110/AEQB [1]));
   XNOR2 \UART_RX_Inst/U89  (.OUT(\UART_RX_Inst/N114 ),
	.B(\UART_RX_Inst/lt_110/AEQB [2]),
	.A(\UART_RX_Inst/n73 ));
   INV \UART_RX_Inst/U88  (.OUT(\UART_RX_Inst/n34 ),
	.IN(\UART_RX_Inst/N184 ));
   INV \UART_RX_Inst/U87  (.OUT(\UART_RX_Inst/n71 ),
	.IN(\UART_RX_Inst/N185 ));
   INV \UART_RX_Inst/U86  (.OUT(\UART_RX_Inst/n72 ),
	.IN(\UART_RX_Inst/r_Clock_Count [0]));
   OAI22 \UART_RX_Inst/U85  (.OUT(\UART_RX_Inst/n165 ),
	.D(\UART_RX_Inst/n72 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n71 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U84  (.OUT(\UART_RX_Inst/n69 ),
	.IN(\UART_RX_Inst/N200 ));
   INV \UART_RX_Inst/U83  (.OUT(\UART_RX_Inst/n70 ),
	.IN(\UART_RX_Inst/r_Clock_Count [15]));
   OAI22 \UART_RX_Inst/U82  (.OUT(\UART_RX_Inst/n164 ),
	.D(\UART_RX_Inst/n70 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n69 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U81  (.OUT(\UART_RX_Inst/n63 ),
	.IN(\UART_RX_Inst/N180 ));
   INV \UART_RX_Inst/U80  (.OUT(\UART_RX_Inst/n67 ),
	.IN(\UART_RX_Inst/N183 ));
   INV \UART_RX_Inst/U79  (.OUT(\UART_RX_Inst/n68 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [2]));
   OAI22 \UART_RX_Inst/U78  (.OUT(\UART_RX_Inst/n163 ),
	.D(\UART_RX_Inst/n68 ),
	.C(\UART_RX_Inst/N180 ),
	.B(\UART_RX_Inst/n67 ),
	.A(\UART_RX_Inst/n63 ));
   INV \UART_RX_Inst/U77  (.OUT(\UART_RX_Inst/n66 ),
	.IN(\UART_RX_Inst/N181 ));
   OAI22 \UART_RX_Inst/U76  (.OUT(\UART_RX_Inst/n162 ),
	.D(\UART_RX_Inst/N112 ),
	.C(\UART_RX_Inst/N180 ),
	.B(\UART_RX_Inst/n66 ),
	.A(\UART_RX_Inst/n63 ));
   INV \UART_RX_Inst/U75  (.OUT(\UART_RX_Inst/n64 ),
	.IN(\UART_RX_Inst/N182 ));
   OAI22 \UART_RX_Inst/U74  (.OUT(\UART_RX_Inst/n161 ),
	.D(\UART_RX_Inst/n65 ),
	.C(\UART_RX_Inst/N180 ),
	.B(\UART_RX_Inst/n64 ),
	.A(\UART_RX_Inst/n63 ));
   INV \UART_RX_Inst/U73  (.OUT(\UART_RX_Inst/n61 ),
	.IN(\UART_RX_Inst/N186 ));
   INV \UART_RX_Inst/U72  (.OUT(\UART_RX_Inst/n62 ),
	.IN(\UART_RX_Inst/r_Clock_Count [1]));
   OAI22 \UART_RX_Inst/U71  (.OUT(\UART_RX_Inst/n160 ),
	.D(\UART_RX_Inst/n62 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n61 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U70  (.OUT(\UART_RX_Inst/n59 ),
	.IN(\UART_RX_Inst/N187 ));
   INV \UART_RX_Inst/U69  (.OUT(\UART_RX_Inst/n60 ),
	.IN(\UART_RX_Inst/r_Clock_Count [2]));
   OAI22 \UART_RX_Inst/U68  (.OUT(\UART_RX_Inst/n159 ),
	.D(\UART_RX_Inst/n60 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n59 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U67  (.OUT(\UART_RX_Inst/n57 ),
	.IN(\UART_RX_Inst/N188 ));
   INV \UART_RX_Inst/U66  (.OUT(\UART_RX_Inst/n58 ),
	.IN(\UART_RX_Inst/r_Clock_Count [3]));
   OAI22 \UART_RX_Inst/U65  (.OUT(\UART_RX_Inst/n158 ),
	.D(\UART_RX_Inst/n58 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n57 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U64  (.OUT(\UART_RX_Inst/n55 ),
	.IN(\UART_RX_Inst/N189 ));
   INV \UART_RX_Inst/U63  (.OUT(\UART_RX_Inst/n56 ),
	.IN(\UART_RX_Inst/r_Clock_Count [4]));
   OAI22 \UART_RX_Inst/U62  (.OUT(\UART_RX_Inst/n157 ),
	.D(\UART_RX_Inst/n56 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n55 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U61  (.OUT(\UART_RX_Inst/n53 ),
	.IN(\UART_RX_Inst/N190 ));
   INV \UART_RX_Inst/U60  (.OUT(\UART_RX_Inst/n54 ),
	.IN(\UART_RX_Inst/r35/AEQB [5]));
   OAI22 \UART_RX_Inst/U59  (.OUT(\UART_RX_Inst/n156 ),
	.D(\UART_RX_Inst/n54 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n53 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U58  (.OUT(\UART_RX_Inst/n51 ),
	.IN(\UART_RX_Inst/N191 ));
   INV \UART_RX_Inst/U57  (.OUT(\UART_RX_Inst/n52 ),
	.IN(\UART_RX_Inst/r_Clock_Count [6]));
   OAI22 \UART_RX_Inst/U56  (.OUT(\UART_RX_Inst/n155 ),
	.D(\UART_RX_Inst/n52 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n51 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U55  (.OUT(\UART_RX_Inst/n49 ),
	.IN(\UART_RX_Inst/N192 ));
   INV \UART_RX_Inst/U54  (.OUT(\UART_RX_Inst/n50 ),
	.IN(\UART_RX_Inst/r_Clock_Count [7]));
   OAI22 \UART_RX_Inst/U53  (.OUT(\UART_RX_Inst/n154 ),
	.D(\UART_RX_Inst/n50 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n49 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U52  (.OUT(\UART_RX_Inst/n47 ),
	.IN(\UART_RX_Inst/N193 ));
   INV \UART_RX_Inst/U51  (.OUT(\UART_RX_Inst/n48 ),
	.IN(\UART_RX_Inst/r35/AEQB [8]));
   OAI22 \UART_RX_Inst/U50  (.OUT(\UART_RX_Inst/n153 ),
	.D(\UART_RX_Inst/n48 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n47 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U49  (.OUT(\UART_RX_Inst/n45 ),
	.IN(\UART_RX_Inst/N194 ));
   INV \UART_RX_Inst/U48  (.OUT(\UART_RX_Inst/n46 ),
	.IN(\UART_RX_Inst/r_Clock_Count [9]));
   OAI22 \UART_RX_Inst/U47  (.OUT(\UART_RX_Inst/n152 ),
	.D(\UART_RX_Inst/n46 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n45 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U46  (.OUT(\UART_RX_Inst/n43 ),
	.IN(\UART_RX_Inst/N195 ));
   INV \UART_RX_Inst/U45  (.OUT(\UART_RX_Inst/n44 ),
	.IN(\UART_RX_Inst/r_Clock_Count [10]));
   OAI22 \UART_RX_Inst/U44  (.OUT(\UART_RX_Inst/n151 ),
	.D(\UART_RX_Inst/n44 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n43 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U43  (.OUT(\UART_RX_Inst/n41 ),
	.IN(\UART_RX_Inst/N196 ));
   INV \UART_RX_Inst/U42  (.OUT(\UART_RX_Inst/n42 ),
	.IN(\UART_RX_Inst/r_Clock_Count [11]));
   OAI22 \UART_RX_Inst/U41  (.OUT(\UART_RX_Inst/n150 ),
	.D(\UART_RX_Inst/n42 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n41 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U40  (.OUT(\UART_RX_Inst/n39 ),
	.IN(\UART_RX_Inst/N197 ));
   INV \UART_RX_Inst/U39  (.OUT(\UART_RX_Inst/n40 ),
	.IN(\UART_RX_Inst/r_Clock_Count [12]));
   OAI22 \UART_RX_Inst/U38  (.OUT(\UART_RX_Inst/n149 ),
	.D(\UART_RX_Inst/n40 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n39 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U37  (.OUT(\UART_RX_Inst/n37 ),
	.IN(\UART_RX_Inst/N198 ));
   INV \UART_RX_Inst/U36  (.OUT(\UART_RX_Inst/n38 ),
	.IN(\UART_RX_Inst/r_Clock_Count [13]));
   OAI22 \UART_RX_Inst/U35  (.OUT(\UART_RX_Inst/n148 ),
	.D(\UART_RX_Inst/n38 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n37 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U34  (.OUT(\UART_RX_Inst/n35 ),
	.IN(\UART_RX_Inst/N199 ));
   INV \UART_RX_Inst/U33  (.OUT(\UART_RX_Inst/n36 ),
	.IN(\UART_RX_Inst/r_Clock_Count [14]));
   OAI22 \UART_RX_Inst/U32  (.OUT(\UART_RX_Inst/n147 ),
	.D(\UART_RX_Inst/n36 ),
	.C(\UART_RX_Inst/N184 ),
	.B(\UART_RX_Inst/n35 ),
	.A(\UART_RX_Inst/n34 ));
   INV \UART_RX_Inst/U31  (.OUT(\UART_RX_Inst/n32 ),
	.IN(\UART_RX_Inst/N201 ));
   INV \UART_RX_Inst/U30  (.OUT(\UART_RX_Inst/n33 ),
	.IN(o_RX_Done));
   OAI22 \UART_RX_Inst/U29  (.OUT(\UART_RX_Inst/n146 ),
	.D(\UART_RX_Inst/n33 ),
	.C(\UART_RX_Inst/N201 ),
	.B(\UART_RX_Inst/n32 ),
	.A(\UART_RX_Inst/n102 ));
   INV \UART_RX_Inst/U28  (.OUT(\UART_RX_Inst/n30 ),
	.IN(\UART_RX_Inst/N213 ));
   INV \UART_RX_Inst/U27  (.OUT(\UART_RX_Inst/n31 ),
	.IN(o_RX_Byte[7]));
   OAI22 \UART_RX_Inst/U26  (.OUT(\UART_RX_Inst/n145 ),
	.D(\UART_RX_Inst/n31 ),
	.C(\UART_RX_Inst/N213 ),
	.B(\UART_RX_Inst/n30 ),
	.A(\UART_RX_Inst/n95 ));
   INV \UART_RX_Inst/U25  (.OUT(\UART_RX_Inst/n28 ),
	.IN(\UART_RX_Inst/N212 ));
   INV \UART_RX_Inst/U24  (.OUT(\UART_RX_Inst/n29 ),
	.IN(o_RX_Byte[6]));
   OAI22 \UART_RX_Inst/U23  (.OUT(\UART_RX_Inst/n144 ),
	.D(\UART_RX_Inst/n29 ),
	.C(\UART_RX_Inst/N212 ),
	.B(\UART_RX_Inst/n28 ),
	.A(\UART_RX_Inst/n95 ));
   INV \UART_RX_Inst/U22  (.OUT(\UART_RX_Inst/n26 ),
	.IN(\UART_RX_Inst/N211 ));
   INV \UART_RX_Inst/U21  (.OUT(\UART_RX_Inst/n27 ),
	.IN(o_RX_Byte[5]));
   OAI22 \UART_RX_Inst/U20  (.OUT(\UART_RX_Inst/n143 ),
	.D(\UART_RX_Inst/n27 ),
	.C(\UART_RX_Inst/N211 ),
	.B(\UART_RX_Inst/n26 ),
	.A(\UART_RX_Inst/n95 ));
   INV \UART_RX_Inst/U19  (.OUT(\UART_RX_Inst/n24 ),
	.IN(\UART_RX_Inst/N210 ));
   INV \UART_RX_Inst/U18  (.OUT(\UART_RX_Inst/n25 ),
	.IN(o_RX_Byte[4]));
   OAI22 \UART_RX_Inst/U17  (.OUT(\UART_RX_Inst/n142 ),
	.D(\UART_RX_Inst/n25 ),
	.C(\UART_RX_Inst/N210 ),
	.B(\UART_RX_Inst/n24 ),
	.A(\UART_RX_Inst/n95 ));
   INV \UART_RX_Inst/U16  (.OUT(\UART_RX_Inst/n22 ),
	.IN(\UART_RX_Inst/N209 ));
   INV \UART_RX_Inst/U15  (.OUT(\UART_RX_Inst/n23 ),
	.IN(o_RX_Byte[3]));
   OAI22 \UART_RX_Inst/U14  (.OUT(\UART_RX_Inst/n141 ),
	.D(\UART_RX_Inst/n23 ),
	.C(\UART_RX_Inst/N209 ),
	.B(\UART_RX_Inst/n22 ),
	.A(\UART_RX_Inst/n95 ));
   INV \UART_RX_Inst/U11  (.OUT(\UART_RX_Inst/n20 ),
	.IN(\UART_RX_Inst/N208 ));
   INV \UART_RX_Inst/U10  (.OUT(\UART_RX_Inst/n21 ),
	.IN(o_RX_Byte[2]));
   OAI22 \UART_RX_Inst/U9  (.OUT(\UART_RX_Inst/n140 ),
	.D(\UART_RX_Inst/n21 ),
	.C(\UART_RX_Inst/N208 ),
	.B(\UART_RX_Inst/n20 ),
	.A(\UART_RX_Inst/n95 ));
   INV \UART_RX_Inst/U8  (.OUT(\UART_RX_Inst/n18 ),
	.IN(\UART_RX_Inst/N207 ));
   INV \UART_RX_Inst/U7  (.OUT(\UART_RX_Inst/n19 ),
	.IN(o_RX_Byte[1]));
   OAI22 \UART_RX_Inst/U6  (.OUT(\UART_RX_Inst/n139 ),
	.D(\UART_RX_Inst/n19 ),
	.C(\UART_RX_Inst/N207 ),
	.B(\UART_RX_Inst/n18 ),
	.A(\UART_RX_Inst/n95 ));
   INV \UART_RX_Inst/U5  (.OUT(\UART_RX_Inst/n16 ),
	.IN(\UART_RX_Inst/N206 ));
   INV \UART_RX_Inst/U4  (.OUT(\UART_RX_Inst/n17 ),
	.IN(o_RX_Byte[0]));
   OAI22 \UART_RX_Inst/U3  (.OUT(\UART_RX_Inst/n138 ),
	.D(\UART_RX_Inst/n17 ),
	.C(\UART_RX_Inst/N206 ),
	.B(\UART_RX_Inst/n16 ),
	.A(\UART_RX_Inst/n95 ));
   DFF \UART_RX_Inst/r_RX_Byte_reg[0]  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Byte[0]),
	.D(\UART_RX_Inst/n138 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_Byte_reg[1]  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Byte[1]),
	.D(\UART_RX_Inst/n139 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_Byte_reg[2]  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Byte[2]),
	.D(\UART_RX_Inst/n140 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_Byte_reg[3]  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Byte[3]),
	.D(\UART_RX_Inst/n141 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_Byte_reg[4]  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Byte[4]),
	.D(\UART_RX_Inst/n142 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_Byte_reg[5]  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Byte[5]),
	.D(\UART_RX_Inst/n143 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_Byte_reg[6]  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Byte[6]),
	.D(\UART_RX_Inst/n144 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_Byte_reg[7]  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Byte[7]),
	.D(\UART_RX_Inst/n145 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[14]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [14]),
	.D(\UART_RX_Inst/n147 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[13]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [13]),
	.D(\UART_RX_Inst/n148 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[12]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [12]),
	.D(\UART_RX_Inst/n149 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[11]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [11]),
	.D(\UART_RX_Inst/n150 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[10]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [10]),
	.D(\UART_RX_Inst/n151 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[9]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [9]),
	.D(\UART_RX_Inst/n152 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[8]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r35/AEQB [8]),
	.D(\UART_RX_Inst/n153 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[7]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [7]),
	.D(\UART_RX_Inst/n154 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[6]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [6]),
	.D(\UART_RX_Inst/n155 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[5]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r35/AEQB [5]),
	.D(\UART_RX_Inst/n156 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[4]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [4]),
	.D(\UART_RX_Inst/n157 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[3]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [3]),
	.D(\UART_RX_Inst/n158 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[2]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [2]),
	.D(\UART_RX_Inst/n159 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[1]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [1]),
	.D(\UART_RX_Inst/n160 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_Done_reg  (.R(\UART_RX_Inst/N21 ),
	.Q(o_RX_Done),
	.D(\UART_RX_Inst/n146 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_State_reg[2]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_RX_State [2]),
	.D(\UART_RX_Inst/N205 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_State_reg[0]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_RX_State [0]),
	.D(\UART_RX_Inst/N203 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Bit_Index_reg[2]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/lt_110/AEQB [2]),
	.D(\UART_RX_Inst/n163 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Bit_Index_reg[1]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/lt_110/AEQB [1]),
	.D(\UART_RX_Inst/n161 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Bit_Index_reg[0]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Bit_Index[0] ),
	.D(\UART_RX_Inst/n162 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_RX_State_reg[1]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_RX_State [1]),
	.D(\UART_RX_Inst/N204 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[15]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [15]),
	.D(\UART_RX_Inst/n164 ),
	.CLK(i_System_Clock));
   DFF \UART_RX_Inst/r_Clock_Count_reg[0]  (.R(\UART_RX_Inst/N21 ),
	.Q(\UART_RX_Inst/r_Clock_Count [0]),
	.D(\UART_RX_Inst/n165 ),
	.CLK(i_System_Clock));
   NAND2 \UART_RX_Inst/C12  (.OUT(\UART_RX_Inst/n83 ),
	.B(\UART_RX_Inst/N24 ),
	.A(\UART_RX_Inst/N23 ));
   NAND2 \UART_RX_Inst/C15  (.OUT(\UART_RX_Inst/N28 ),
	.B(\UART_RX_Inst/N24 ),
	.A(\UART_RX_Inst/N23 ));
   NAND2 \UART_RX_Inst/C19  (.OUT(\UART_RX_Inst/N31 ),
	.B(\UART_RX_Inst/r_RX_State [1]),
	.A(\UART_RX_Inst/N23 ));
   NAND2 \UART_RX_Inst/C24  (.OUT(\UART_RX_Inst/N34 ),
	.B(\UART_RX_Inst/r_RX_State [1]),
	.A(\UART_RX_Inst/N23 ));
   NAND2 \UART_RX_Inst/C28  (.OUT(\UART_RX_Inst/N37 ),
	.B(\UART_RX_Inst/N24 ),
	.A(\UART_RX_Inst/r_RX_State [2]));
   NAND2 \UART_RX_Inst/C320  (.OUT(\UART_RX_Inst/n130 ),
	.B(\UART_RX_Inst/lt_110/AEQB [1]),
	.A(\UART_RX_Inst/r_Bit_Index[0] ));
   NAND2 \UART_RX_Inst/C321  (.OUT(\UART_RX_Inst/n82 ),
	.B(\UART_RX_Inst/lt_110/AEQB [2]),
	.A(\UART_RX_Inst/N219 ));
   NAND2 \UART_RX_Inst/C322  (.OUT(\UART_RX_Inst/n131 ),
	.B(\UART_RX_Inst/lt_110/AEQB [1]),
	.A(\UART_RX_Inst/N0 ));
   INV \UART_RX_Inst/I_1  (.OUT(\UART_RX_Inst/N0 ),
	.IN(\UART_RX_Inst/r_Bit_Index[0] ));
   NAND2 \UART_RX_Inst/C323  (.OUT(\UART_RX_Inst/n81 ),
	.B(\UART_RX_Inst/lt_110/AEQB [2]),
	.A(\UART_RX_Inst/N220 ));
   NAND2 \UART_RX_Inst/C324  (.OUT(\UART_RX_Inst/n132 ),
	.B(\UART_RX_Inst/N1 ),
	.A(\UART_RX_Inst/r_Bit_Index[0] ));
   INV \UART_RX_Inst/I_2  (.OUT(\UART_RX_Inst/N1 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [1]));
   NAND2 \UART_RX_Inst/C325  (.OUT(\UART_RX_Inst/n80 ),
	.B(\UART_RX_Inst/lt_110/AEQB [2]),
	.A(\UART_RX_Inst/N221 ));
   NAND2 \UART_RX_Inst/C326  (.OUT(\UART_RX_Inst/n133 ),
	.B(\UART_RX_Inst/N3 ),
	.A(\UART_RX_Inst/N2 ));
   INV \UART_RX_Inst/I_3  (.OUT(\UART_RX_Inst/N2 ),
	.IN(\UART_RX_Inst/r_Bit_Index[0] ));
   INV \UART_RX_Inst/I_4  (.OUT(\UART_RX_Inst/N3 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [1]));
   NAND2 \UART_RX_Inst/C327  (.OUT(\UART_RX_Inst/n79 ),
	.B(\UART_RX_Inst/lt_110/AEQB [2]),
	.A(\UART_RX_Inst/N222 ));
   NAND2 \UART_RX_Inst/C328  (.OUT(\UART_RX_Inst/n134 ),
	.B(\UART_RX_Inst/lt_110/AEQB [1]),
	.A(\UART_RX_Inst/r_Bit_Index[0] ));
   NAND2 \UART_RX_Inst/C329  (.OUT(\UART_RX_Inst/n78 ),
	.B(\UART_RX_Inst/N4 ),
	.A(\UART_RX_Inst/N223 ));
   INV \UART_RX_Inst/I_5  (.OUT(\UART_RX_Inst/N4 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [2]));
   NAND2 \UART_RX_Inst/C330  (.OUT(\UART_RX_Inst/n135 ),
	.B(\UART_RX_Inst/lt_110/AEQB [1]),
	.A(\UART_RX_Inst/N5 ));
   INV \UART_RX_Inst/I_6  (.OUT(\UART_RX_Inst/N5 ),
	.IN(\UART_RX_Inst/r_Bit_Index[0] ));
   NAND2 \UART_RX_Inst/C331  (.OUT(\UART_RX_Inst/n77 ),
	.B(\UART_RX_Inst/N6 ),
	.A(\UART_RX_Inst/N224 ));
   INV \UART_RX_Inst/I_7  (.OUT(\UART_RX_Inst/N6 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [2]));
   NAND2 \UART_RX_Inst/C332  (.OUT(\UART_RX_Inst/n136 ),
	.B(\UART_RX_Inst/N7 ),
	.A(\UART_RX_Inst/r_Bit_Index[0] ));
   INV \UART_RX_Inst/I_8  (.OUT(\UART_RX_Inst/N7 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [1]));
   NAND2 \UART_RX_Inst/C333  (.OUT(\UART_RX_Inst/n76 ),
	.B(\UART_RX_Inst/N8 ),
	.A(\UART_RX_Inst/N225 ));
   INV \UART_RX_Inst/I_9  (.OUT(\UART_RX_Inst/N8 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [2]));
   NAND2 \UART_RX_Inst/C334  (.OUT(\UART_RX_Inst/n137 ),
	.B(\UART_RX_Inst/N10 ),
	.A(\UART_RX_Inst/N9 ));
   INV \UART_RX_Inst/I_10  (.OUT(\UART_RX_Inst/N9 ),
	.IN(\UART_RX_Inst/r_Bit_Index[0] ));
   INV \UART_RX_Inst/I_11  (.OUT(\UART_RX_Inst/N10 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [1]));
   NAND2 \UART_RX_Inst/C335  (.OUT(\UART_RX_Inst/n75 ),
	.B(\UART_RX_Inst/N11 ),
	.A(\UART_RX_Inst/N226 ));
   INV \UART_RX_Inst/I_12  (.OUT(\UART_RX_Inst/N11 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [2]));
   INV \UART_RX_Inst/I_14  (.OUT(\UART_RX_Inst/N21 ),
	.IN(i_Rst_L));
   INV \UART_RX_Inst/I_15  (.OUT(\UART_RX_Inst/N23 ),
	.IN(\UART_RX_Inst/r_RX_State [2]));
   INV \UART_RX_Inst/I_16  (.OUT(\UART_RX_Inst/N24 ),
	.IN(\UART_RX_Inst/r_RX_State [1]));
   INV \UART_RX_Inst/I_18  (.OUT(\UART_RX_Inst/U3/U1/Z_7 ),
	.IN(\UART_RX_Inst/N29 ));
   INV \UART_RX_Inst/I_19  (.OUT(\UART_RX_Inst/N33 ),
	.IN(\UART_RX_Inst/N32 ));
   INV \UART_RX_Inst/I_20  (.OUT(\UART_RX_Inst/N202 ),
	.IN(\UART_RX_Inst/N35 ));
   INV \UART_RX_Inst/I_21  (.OUT(\UART_RX_Inst/N39 ),
	.IN(\UART_RX_Inst/N38 ));
   NAND2 \UART_RX_Inst/lt_110/ULTI2  (.OUT(\UART_RX_Inst/N84 ),
	.B(\UART_RX_Inst/lt_110/LTV2 [2]),
	.A(\UART_RX_Inst/lt_110/LTV1 [2]));
   NAND2 \UART_RX_Inst/lt_110/ULTI1  (.OUT(\UART_RX_Inst/lt_110/LTV2 [2]),
	.B(\UART_RX_Inst/lt_110/LTV [2]),
	.A(\UART_RX_Inst/lt_110/AEQB [2]));
   NAND2 \UART_RX_Inst/lt_110/ULTI2_1  (.OUT(\UART_RX_Inst/lt_110/LTV [2]),
	.B(\UART_RX_Inst/lt_110/LTV2 [1]),
	.A(\UART_RX_Inst/lt_110/LTV1 [1]));
   NAND2 \UART_RX_Inst/lt_110/ULTI1_1  (.OUT(\UART_RX_Inst/lt_110/LTV2 [1]),
	.B(\UART_RX_Inst/lt_110/LTV [1]),
	.A(\UART_RX_Inst/lt_110/AEQB [1]));
   OAI22 \UART_TX_Inst/U147  (.OUT(\UART_TX_Inst/n122 ),
	.D(\UART_TX_Inst/n119 ),
	.C(\UART_TX_Inst/lt_109/AEQB [1]),
	.B(\UART_TX_Inst/n121 ),
	.A(\UART_TX_Inst/n108 ));
   INV \UART_TX_Inst/U146  (.OUT(\UART_TX_Inst/n121 ),
	.IN(\UART_TX_Inst/n120 ));
   OAI22 \UART_TX_Inst/U145  (.OUT(\UART_TX_Inst/n120 ),
	.D(\UART_TX_Inst/n111 ),
	.C(\UART_TX_Inst/N9 ),
	.B(\UART_TX_Inst/n112 ),
	.A(\UART_TX_Inst/n104 ));
   INV \UART_TX_Inst/U144  (.OUT(\UART_TX_Inst/n119 ),
	.IN(\UART_TX_Inst/n118 ));
   OAI22 \UART_TX_Inst/U143  (.OUT(\UART_TX_Inst/n118 ),
	.D(\UART_TX_Inst/n109 ),
	.C(\UART_TX_Inst/N9 ),
	.B(\UART_TX_Inst/n110 ),
	.A(\UART_TX_Inst/n104 ));
   OAI22 \UART_TX_Inst/U142  (.OUT(\UART_TX_Inst/n117 ),
	.D(\UART_TX_Inst/n114 ),
	.C(\UART_TX_Inst/lt_109/AEQB [1]),
	.B(\UART_TX_Inst/n108 ),
	.A(\UART_TX_Inst/n116 ));
   INV \UART_TX_Inst/U141  (.OUT(\UART_TX_Inst/n116 ),
	.IN(\UART_TX_Inst/n115 ));
   OAI22 \UART_TX_Inst/U140  (.OUT(\UART_TX_Inst/n115 ),
	.D(\UART_TX_Inst/n106 ),
	.C(\UART_TX_Inst/N9 ),
	.B(\UART_TX_Inst/n107 ),
	.A(\UART_TX_Inst/n104 ));
   INV \UART_TX_Inst/U139  (.OUT(\UART_TX_Inst/n114 ),
	.IN(\UART_TX_Inst/n113 ));
   OAI22 \UART_TX_Inst/U138  (.OUT(\UART_TX_Inst/n113 ),
	.D(\UART_TX_Inst/n103 ),
	.C(\UART_TX_Inst/N9 ),
	.B(\UART_TX_Inst/n105 ),
	.A(\UART_TX_Inst/n104 ));
   INV \UART_TX_Inst/U137  (.OUT(\UART_TX_Inst/n112 ),
	.IN(\UART_TX_Inst/r_TX_Data [7]));
   INV \UART_TX_Inst/U136  (.OUT(\UART_TX_Inst/n111 ),
	.IN(\UART_TX_Inst/r_TX_Data [6]));
   INV \UART_TX_Inst/U135  (.OUT(\UART_TX_Inst/n110 ),
	.IN(\UART_TX_Inst/r_TX_Data [5]));
   INV \UART_TX_Inst/U134  (.OUT(\UART_TX_Inst/n109 ),
	.IN(\UART_TX_Inst/r_TX_Data [4]));
   INV \UART_TX_Inst/U133  (.OUT(\UART_TX_Inst/n108 ),
	.IN(\UART_TX_Inst/lt_109/AEQB [1]));
   INV \UART_TX_Inst/U132  (.OUT(\UART_TX_Inst/n107 ),
	.IN(\UART_TX_Inst/r_TX_Data [3]));
   INV \UART_TX_Inst/U131  (.OUT(\UART_TX_Inst/n106 ),
	.IN(\UART_TX_Inst/r_TX_Data [2]));
   INV \UART_TX_Inst/U130  (.OUT(\UART_TX_Inst/n105 ),
	.IN(\UART_TX_Inst/r_TX_Data [1]));
   INV \UART_TX_Inst/U129  (.OUT(\UART_TX_Inst/n104 ),
	.IN(\UART_TX_Inst/N9 ));
   INV \UART_TX_Inst/U128  (.OUT(\UART_TX_Inst/n103 ),
	.IN(\UART_TX_Inst/r_TX_Data [0]));
   INV \UART_TX_Inst/U127  (.OUT(\UART_TX_Inst/N66 ),
	.IN(\UART_TX_Inst/N9 ));
   INV \UART_TX_Inst/U126  (.OUT(\UART_TX_Inst/n102 ),
	.IN(\UART_TX_Inst/lt_109/AEQB [1]));
   INV \UART_TX_Inst/U121  (.OUT(\UART_TX_Inst/n88 ),
	.IN(\UART_TX_Inst/N144 ));
   INV \UART_TX_Inst/U120  (.OUT(\UART_TX_Inst/n87 ),
	.IN(\UART_TX_Inst/N143 ));
   INV \UART_TX_Inst/U119  (.OUT(\UART_TX_Inst/n86 ),
	.IN(\UART_TX_Inst/N142 ));
   INV \UART_TX_Inst/U118  (.OUT(\UART_TX_Inst/n85 ),
	.IN(\UART_TX_Inst/r_Clock_Count [2]));
   INV \UART_TX_Inst/U117  (.OUT(\UART_TX_Inst/n84 ),
	.IN(\UART_TX_Inst/N141 ));
   INV \UART_TX_Inst/U116  (.OUT(\UART_TX_Inst/n83 ),
	.IN(\UART_TX_Inst/r_Clock_Count [3]));
   INV \UART_TX_Inst/U115  (.OUT(\UART_TX_Inst/n82 ),
	.IN(\UART_TX_Inst/N140 ));
   INV \UART_TX_Inst/U114  (.OUT(\UART_TX_Inst/n81 ),
	.IN(\UART_TX_Inst/r_Clock_Count [4]));
   INV \UART_TX_Inst/U113  (.OUT(\UART_TX_Inst/n80 ),
	.IN(\UART_TX_Inst/N139 ));
   INV \UART_TX_Inst/U112  (.OUT(\UART_TX_Inst/n79 ),
	.IN(\UART_TX_Inst/N138 ));
   INV \UART_TX_Inst/U111  (.OUT(\UART_TX_Inst/n78 ),
	.IN(\UART_TX_Inst/N137 ));
   INV \UART_TX_Inst/U110  (.OUT(\UART_TX_Inst/n77 ),
	.IN(\UART_TX_Inst/r_Clock_Count [7]));
   INV \UART_TX_Inst/U109  (.OUT(\UART_TX_Inst/n76 ),
	.IN(\UART_TX_Inst/N136 ));
   INV \UART_TX_Inst/U108  (.OUT(\UART_TX_Inst/n75 ),
	.IN(\UART_TX_Inst/r_Clock_Count [10]));
   INV \UART_TX_Inst/U107  (.OUT(\UART_TX_Inst/n74 ),
	.IN(\UART_TX_Inst/N18 ));
   INV \UART_TX_Inst/U106  (.OUT(\UART_TX_Inst/n48 ),
	.IN(\UART_TX_Inst/N23 ));
   OAI22 \UART_TX_Inst/U105  (.OUT(\UART_TX_Inst/n53 ),
	.D(\UART_TX_Inst/n50 ),
	.C(\UART_TX_Inst/N146 ),
	.B(\UART_TX_Inst/n48 ),
	.A(\UART_TX_Inst/n74 ));
   INV \UART_TX_Inst/U104  (.OUT(\UART_TX_Inst/n46 ),
	.IN(\UART_TX_Inst/N20 ));
   NOR2 \UART_TX_Inst/U103  (.OUT(\UART_TX_Inst/n73 ),
	.B(\UART_TX_Inst/n48 ),
	.A(\UART_TX_Inst/n46 ));
   NOR2 \UART_TX_Inst/U102  (.OUT(\UART_TX_Inst/n61 ),
	.B(\UART_TX_Inst/n73 ),
	.A(\UART_TX_Inst/n53 ));
   INV \UART_TX_Inst/U101  (.OUT(\UART_TX_Inst/n72 ),
	.IN(\UART_TX_Inst/N87 ));
   NOR2 \UART_TX_Inst/U100  (.OUT(\UART_TX_Inst/N110 ),
	.B(\UART_TX_Inst/n72 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U99  (.OUT(\UART_TX_Inst/n71 ),
	.IN(\UART_TX_Inst/N88 ));
   NOR2 \UART_TX_Inst/U98  (.OUT(\UART_TX_Inst/N111 ),
	.B(\UART_TX_Inst/n71 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U97  (.OUT(\UART_TX_Inst/n70 ),
	.IN(\UART_TX_Inst/N89 ));
   NOR2 \UART_TX_Inst/U96  (.OUT(\UART_TX_Inst/N112 ),
	.B(\UART_TX_Inst/n70 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U95  (.OUT(\UART_TX_Inst/n69 ),
	.IN(\UART_TX_Inst/N90 ));
   NOR2 \UART_TX_Inst/U94  (.OUT(\UART_TX_Inst/N113 ),
	.B(\UART_TX_Inst/n69 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U93  (.OUT(\UART_TX_Inst/n68 ),
	.IN(\UART_TX_Inst/N91 ));
   NOR2 \UART_TX_Inst/U92  (.OUT(\UART_TX_Inst/N114 ),
	.B(\UART_TX_Inst/n68 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U91  (.OUT(\UART_TX_Inst/n67 ),
	.IN(\UART_TX_Inst/N92 ));
   NOR2 \UART_TX_Inst/U90  (.OUT(\UART_TX_Inst/N115 ),
	.B(\UART_TX_Inst/n67 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U89  (.OUT(\UART_TX_Inst/n66 ),
	.IN(\UART_TX_Inst/N93 ));
   NOR2 \UART_TX_Inst/U88  (.OUT(\UART_TX_Inst/N116 ),
	.B(\UART_TX_Inst/n66 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U87  (.OUT(\UART_TX_Inst/n65 ),
	.IN(\UART_TX_Inst/N94 ));
   NOR2 \UART_TX_Inst/U86  (.OUT(\UART_TX_Inst/N117 ),
	.B(\UART_TX_Inst/n65 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U85  (.OUT(\UART_TX_Inst/n64 ),
	.IN(\UART_TX_Inst/N95 ));
   NOR2 \UART_TX_Inst/U84  (.OUT(\UART_TX_Inst/N118 ),
	.B(\UART_TX_Inst/n64 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U83  (.OUT(\UART_TX_Inst/n63 ),
	.IN(\UART_TX_Inst/N96 ));
   NOR2 \UART_TX_Inst/U82  (.OUT(\UART_TX_Inst/N119 ),
	.B(\UART_TX_Inst/n63 ),
	.A(\UART_TX_Inst/n61 ));
   INV \UART_TX_Inst/U81  (.OUT(\UART_TX_Inst/n62 ),
	.IN(\UART_TX_Inst/N97 ));
   NOR2 \UART_TX_Inst/U80  (.OUT(\UART_TX_Inst/N120 ),
	.B(\UART_TX_Inst/n62 ),
	.A(\UART_TX_Inst/n61 ));
   NAND2 \UART_TX_Inst/U79  (.OUT(\UART_TX_Inst/n60 ),
	.B(\UART_TX_Inst/n48 ),
	.A(\UART_TX_Inst/N20 ));
   NAND2 \UART_TX_Inst/U78  (.OUT(\UART_TX_Inst/N121 ),
	.B(\UART_TX_Inst/n60 ),
	.A(\UART_TX_Inst/n59 ));
   NAND2 \UART_TX_Inst/U77  (.OUT(\UART_TX_Inst/n55 ),
	.B(\UART_TX_Inst/N20 ),
	.A(\UART_TX_Inst/N64 ));
   INV \UART_TX_Inst/U76  (.OUT(\UART_TX_Inst/n58 ),
	.IN(\UART_TX_Inst/N66 ));
   NOR2 \UART_TX_Inst/U75  (.OUT(\UART_TX_Inst/N122 ),
	.B(\UART_TX_Inst/n58 ),
	.A(\UART_TX_Inst/n55 ));
   INV \UART_TX_Inst/U74  (.OUT(\UART_TX_Inst/n57 ),
	.IN(\UART_TX_Inst/N67 ));
   NOR2 \UART_TX_Inst/U73  (.OUT(\UART_TX_Inst/N123 ),
	.B(\UART_TX_Inst/n57 ),
	.A(\UART_TX_Inst/n55 ));
   INV \UART_TX_Inst/U72  (.OUT(\UART_TX_Inst/n56 ),
	.IN(\UART_TX_Inst/N68 ));
   NOR2 \UART_TX_Inst/U71  (.OUT(\UART_TX_Inst/N124 ),
	.B(\UART_TX_Inst/n56 ),
	.A(\UART_TX_Inst/n55 ));
   INV \UART_TX_Inst/U70  (.OUT(\UART_TX_Inst/n54 ),
	.IN(\UART_TX_Inst/N64 ));
   NAND3 \UART_TX_Inst/U69  (.OUT(\UART_TX_Inst/n51 ),
	.C(\UART_TX_Inst/N20 ),
	.B(\UART_TX_Inst/n54 ),
	.A(\UART_TX_Inst/n48 ));
   NAND2 \UART_TX_Inst/U68  (.OUT(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/N16 ),
	.A(i_TX_Valid));
   INV \UART_TX_Inst/U67  (.OUT(\UART_TX_Inst/n52 ),
	.IN(\UART_TX_Inst/n53 ));
   NAND3 \UART_TX_Inst/U66  (.OUT(\UART_TX_Inst/N125 ),
	.C(\UART_TX_Inst/n52 ),
	.B(\UART_TX_Inst/n43 ),
	.A(\UART_TX_Inst/n51 ));
   INV \UART_TX_Inst/U65  (.OUT(\UART_TX_Inst/n44 ),
	.IN(\UART_TX_Inst/n50 ));
   INV \UART_TX_Inst/U64  (.OUT(\UART_TX_Inst/n49 ),
	.IN(\UART_TX_Inst/N146 ));
   NAND2 \UART_TX_Inst/U63  (.OUT(\UART_TX_Inst/n45 ),
	.B(\UART_TX_Inst/n49 ),
	.A(\UART_TX_Inst/n44 ));
   NAND2 \UART_TX_Inst/U62  (.OUT(\UART_TX_Inst/n47 ),
	.B(\UART_TX_Inst/n48 ),
	.A(\UART_TX_Inst/N18 ));
   NAND3 \UART_TX_Inst/U61  (.OUT(\UART_TX_Inst/N126 ),
	.C(\UART_TX_Inst/n47 ),
	.B(\UART_TX_Inst/n46 ),
	.A(\UART_TX_Inst/n45 ));
   NAND2 \UART_TX_Inst/U60  (.OUT(\UART_TX_Inst/n42 ),
	.B(\UART_TX_Inst/n44 ),
	.A(\UART_TX_Inst/N146 ));
   NAND2 \UART_TX_Inst/U59  (.OUT(\UART_TX_Inst/N127 ),
	.B(\UART_TX_Inst/n43 ),
	.A(\UART_TX_Inst/n42 ));
   INV \UART_TX_Inst/U58  (.OUT(\UART_TX_Inst/N129 ),
	.IN(\UART_TX_Inst/n42 ));
   INV \UART_TX_Inst/U57  (.OUT(\UART_TX_Inst/n41 ),
	.IN(\UART_TX_Inst/r_SM_Main [1]));
   NAND2 \UART_TX_Inst/U56  (.OUT(\UART_TX_Inst/N17 ),
	.B(\UART_TX_Inst/n41 ),
	.A(\UART_TX_Inst/r_SM_Main [0]));
   INV \UART_TX_Inst/U53  (.OUT(\UART_TX_Inst/n37 ),
	.IN(\UART_TX_Inst/r_SM_Main [1]));
   NOR2 \UART_TX_Inst/U52  (.OUT(\UART_TX_Inst/N20 ),
	.B(\UART_TX_Inst/r_SM_Main [0]),
	.A(\UART_TX_Inst/n37 ));
   NAND2 \UART_TX_Inst/U51  (.OUT(\UART_TX_Inst/n36 ),
	.B(\UART_TX_Inst/n37 ),
	.A(\UART_TX_Inst/r_SM_Main [0]));
   INV \UART_TX_Inst/U50  (.OUT(\UART_TX_Inst/n35 ),
	.IN(\UART_TX_Inst/n36 ));
   NOR2 \UART_TX_Inst/U49  (.OUT(\UART_TX_Inst/n11 ),
	.B(\UART_TX_Inst/n35 ),
	.A(\UART_TX_Inst/N20 ));
   NAND2 \UART_TX_Inst/U48  (.OUT(\UART_TX_Inst/n50 ),
	.B(\UART_TX_Inst/r_SM_Main [1]),
	.A(\UART_TX_Inst/r_SM_Main [0]));
   NAND2 \UART_TX_Inst/U47  (.OUT(\UART_TX_Inst/n59 ),
	.B(\UART_TX_Inst/n50 ),
	.A(\UART_TX_Inst/n11 ));
   INV \UART_TX_Inst/U46  (.OUT(\UART_TX_Inst/N16 ),
	.IN(\UART_TX_Inst/n59 ));
   XNOR2 \UART_TX_Inst/U45  (.OUT(\UART_TX_Inst/n34 ),
	.B(\UART_TX_Inst/N66 ),
	.A(\UART_TX_Inst/n102 ));
   INV \UART_TX_Inst/U44  (.OUT(\UART_TX_Inst/N67 ),
	.IN(\UART_TX_Inst/n34 ));
   INV \UART_TX_Inst/U43  (.OUT(\UART_TX_Inst/n15 ),
	.IN(\UART_TX_Inst/lt_109/AEQB [2]));
   NOR2 \UART_TX_Inst/U42  (.OUT(\UART_TX_Inst/n33 ),
	.B(\UART_TX_Inst/N66 ),
	.A(\UART_TX_Inst/n102 ));
   XNOR2 \UART_TX_Inst/U41  (.OUT(\UART_TX_Inst/N68 ),
	.B(\UART_TX_Inst/n33 ),
	.A(\UART_TX_Inst/n15 ));
   INV \UART_TX_Inst/U40  (.OUT(\UART_TX_Inst/n29 ),
	.IN(\UART_TX_Inst/N121 ));
   INV \UART_TX_Inst/U39  (.OUT(\UART_TX_Inst/n32 ),
	.IN(\UART_TX_Inst/N124 ));
   OAI22 \UART_TX_Inst/U38  (.OUT(\UART_TX_Inst/n100 ),
	.D(\UART_TX_Inst/n15 ),
	.C(\UART_TX_Inst/N121 ),
	.B(\UART_TX_Inst/n32 ),
	.A(\UART_TX_Inst/n29 ));
   INV \UART_TX_Inst/U37  (.OUT(\UART_TX_Inst/n31 ),
	.IN(\UART_TX_Inst/N122 ));
   OAI22 \UART_TX_Inst/U36  (.OUT(\UART_TX_Inst/n99 ),
	.D(\UART_TX_Inst/N121 ),
	.C(\UART_TX_Inst/N66 ),
	.B(\UART_TX_Inst/n31 ),
	.A(\UART_TX_Inst/n29 ));
   INV \UART_TX_Inst/U35  (.OUT(\UART_TX_Inst/n30 ),
	.IN(\UART_TX_Inst/N123 ));
   OAI22 \UART_TX_Inst/U34  (.OUT(\UART_TX_Inst/n98 ),
	.D(\UART_TX_Inst/N121 ),
	.C(\UART_TX_Inst/n102 ),
	.B(\UART_TX_Inst/n30 ),
	.A(\UART_TX_Inst/n29 ));
   INV \UART_TX_Inst/U33  (.OUT(\UART_TX_Inst/n27 ),
	.IN(\UART_TX_Inst/N127 ));
   INV \UART_TX_Inst/U32  (.OUT(\UART_TX_Inst/n28 ),
	.IN(o_TX_Busy));
   OAI22 \UART_TX_Inst/U31  (.OUT(\UART_TX_Inst/n97 ),
	.D(\UART_TX_Inst/n28 ),
	.C(\UART_TX_Inst/N127 ),
	.B(\UART_TX_Inst/n27 ),
	.A(\UART_TX_Inst/n59 ));
   INV \UART_TX_Inst/U30  (.OUT(\UART_TX_Inst/n18 ),
	.IN(\UART_TX_Inst/n43 ));
   INV \UART_TX_Inst/U29  (.OUT(\UART_TX_Inst/n26 ),
	.IN(i_TX_Byte[0]));
   OAI22 \UART_TX_Inst/U28  (.OUT(\UART_TX_Inst/n96 ),
	.D(\UART_TX_Inst/n26 ),
	.C(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/n103 ),
	.A(\UART_TX_Inst/n18 ));
   INV \UART_TX_Inst/U27  (.OUT(\UART_TX_Inst/n25 ),
	.IN(i_TX_Byte[1]));
   OAI22 \UART_TX_Inst/U26  (.OUT(\UART_TX_Inst/n95 ),
	.D(\UART_TX_Inst/n25 ),
	.C(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/n105 ),
	.A(\UART_TX_Inst/n18 ));
   INV \UART_TX_Inst/U25  (.OUT(\UART_TX_Inst/n24 ),
	.IN(i_TX_Byte[2]));
   OAI22 \UART_TX_Inst/U24  (.OUT(\UART_TX_Inst/n94 ),
	.D(\UART_TX_Inst/n24 ),
	.C(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/n106 ),
	.A(\UART_TX_Inst/n18 ));
   INV \UART_TX_Inst/U23  (.OUT(\UART_TX_Inst/n23 ),
	.IN(i_TX_Byte[3]));
   OAI22 \UART_TX_Inst/U22  (.OUT(\UART_TX_Inst/n93 ),
	.D(\UART_TX_Inst/n23 ),
	.C(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/n107 ),
	.A(\UART_TX_Inst/n18 ));
   INV \UART_TX_Inst/U21  (.OUT(\UART_TX_Inst/n22 ),
	.IN(i_TX_Byte[4]));
   OAI22 \UART_TX_Inst/U20  (.OUT(\UART_TX_Inst/n92 ),
	.D(\UART_TX_Inst/n22 ),
	.C(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/n109 ),
	.A(\UART_TX_Inst/n18 ));
   INV \UART_TX_Inst/U19  (.OUT(\UART_TX_Inst/n21 ),
	.IN(i_TX_Byte[5]));
   OAI22 \UART_TX_Inst/U18  (.OUT(\UART_TX_Inst/n91 ),
	.D(\UART_TX_Inst/n21 ),
	.C(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/n110 ),
	.A(\UART_TX_Inst/n18 ));
   INV \UART_TX_Inst/U17  (.OUT(\UART_TX_Inst/n20 ),
	.IN(i_TX_Byte[6]));
   OAI22 \UART_TX_Inst/U16  (.OUT(\UART_TX_Inst/n90 ),
	.D(\UART_TX_Inst/n20 ),
	.C(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/n111 ),
	.A(\UART_TX_Inst/n18 ));
   INV \UART_TX_Inst/U15  (.OUT(\UART_TX_Inst/n19 ),
	.IN(i_TX_Byte[7]));
   OAI22 \UART_TX_Inst/U14  (.OUT(\UART_TX_Inst/n89 ),
	.D(\UART_TX_Inst/n19 ),
	.C(\UART_TX_Inst/n43 ),
	.B(\UART_TX_Inst/n112 ),
	.A(\UART_TX_Inst/n18 ));
   INV \UART_TX_Inst/U13  (.OUT(\UART_TX_Inst/n8 ),
	.IN(o_TX_Serial));
   INV \UART_TX_Inst/U10  (.OUT(\UART_TX_Inst/n16 ),
	.IN(\UART_TX_Inst/n122 ));
   INV \UART_TX_Inst/U9  (.OUT(\UART_TX_Inst/n17 ),
	.IN(\UART_TX_Inst/n117 ));
   OAI22 \UART_TX_Inst/U8  (.OUT(\UART_TX_Inst/n14 ),
	.D(\UART_TX_Inst/n17 ),
	.C(\UART_TX_Inst/lt_109/AEQB [2]),
	.B(\UART_TX_Inst/n16 ),
	.A(\UART_TX_Inst/n15 ));
   NAND2 \UART_TX_Inst/U7  (.OUT(\UART_TX_Inst/n13 ),
	.B(\UART_TX_Inst/n14 ),
	.A(\UART_TX_Inst/r_SM_Main [1]));
   INV \UART_TX_Inst/U6  (.OUT(\UART_TX_Inst/n12 ),
	.IN(\UART_TX_Inst/n13 ));
   NOR2 \UART_TX_Inst/U5  (.OUT(\UART_TX_Inst/n9 ),
	.B(\UART_TX_Inst/n12 ),
	.A(\UART_TX_Inst/n11 ));
   INV \UART_TX_Inst/U4  (.OUT(\UART_TX_Inst/n10 ),
	.IN(i_Rst_L));
   OAI22 \UART_TX_Inst/U3  (.OUT(\UART_TX_Inst/n39 ),
	.D(\UART_TX_Inst/n10 ),
	.C(\UART_TX_Inst/n9 ),
	.B(\UART_TX_Inst/n8 ),
	.A(i_Rst_L));
   DFF \UART_TX_Inst/o_TX_Serial_reg  (.R(1'b0),
	.Q(o_TX_Serial),
	.D(\UART_TX_Inst/n39 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Bit_Index_reg[2]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/lt_109/AEQB [2]),
	.D(\UART_TX_Inst/n100 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Bit_Index_reg[1]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/lt_109/AEQB [1]),
	.D(\UART_TX_Inst/n98 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Bit_Index_reg[0]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/N9 ),
	.D(\UART_TX_Inst/n99 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/o_TX_Busy_reg  (.R(\UART_TX_Inst/N12 ),
	.Q(o_TX_Busy),
	.D(\UART_TX_Inst/n97 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/o_TX_Done_reg  (.R(\UART_TX_Inst/N12 ),
	.Q(o_TX_Done),
	.D(\UART_TX_Inst/N129 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_TX_Data_reg[7]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_TX_Data [7]),
	.D(\UART_TX_Inst/n89 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_TX_Data_reg[6]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_TX_Data [6]),
	.D(\UART_TX_Inst/n90 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_TX_Data_reg[5]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_TX_Data [5]),
	.D(\UART_TX_Inst/n91 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_TX_Data_reg[4]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_TX_Data [4]),
	.D(\UART_TX_Inst/n92 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_TX_Data_reg[3]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_TX_Data [3]),
	.D(\UART_TX_Inst/n93 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_TX_Data_reg[2]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_TX_Data [2]),
	.D(\UART_TX_Inst/n94 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_TX_Data_reg[1]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_TX_Data [1]),
	.D(\UART_TX_Inst/n95 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_TX_Data_reg[0]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_TX_Data [0]),
	.D(\UART_TX_Inst/n96 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_SM_Main_reg[1]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_SM_Main [1]),
	.D(\UART_TX_Inst/N126 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[10]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_Clock_Count [10]),
	.D(\UART_TX_Inst/N120 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[9]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r31/AEQB [9]),
	.D(\UART_TX_Inst/N119 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[8]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r31/AEQB [8]),
	.D(\UART_TX_Inst/N118 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[7]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_Clock_Count [7]),
	.D(\UART_TX_Inst/N117 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[6]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r31/AEQB [6]),
	.D(\UART_TX_Inst/N116 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[5]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r31/AEQB [5]),
	.D(\UART_TX_Inst/N115 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[4]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_Clock_Count [4]),
	.D(\UART_TX_Inst/N114 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[3]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_Clock_Count [3]),
	.D(\UART_TX_Inst/N113 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[2]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_Clock_Count [2]),
	.D(\UART_TX_Inst/N112 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[1]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r31/AEQB [1]),
	.D(\UART_TX_Inst/N111 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_Clock_Count_reg[0]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_Clock_Count [0]),
	.D(\UART_TX_Inst/N110 ),
	.CLK(i_System_Clock));
   DFF \UART_TX_Inst/r_SM_Main_reg[0]  (.R(\UART_TX_Inst/N12 ),
	.Q(\UART_TX_Inst/r_SM_Main [0]),
	.D(\UART_TX_Inst/N125 ),
	.CLK(i_System_Clock));
   NAND2 \UART_TX_Inst/C222  (.OUT(\UART_TX_Inst/N136 ),
	.B(\UART_TX_Inst/n75 ),
	.A(\UART_TX_Inst/r31/AEQB [9]));
   NAND2 \UART_TX_Inst/C223  (.OUT(\UART_TX_Inst/N137 ),
	.B(\UART_TX_Inst/n76 ),
	.A(\UART_TX_Inst/r31/AEQB [8]));
   NAND2 \UART_TX_Inst/C224  (.OUT(\UART_TX_Inst/N138 ),
	.B(\UART_TX_Inst/n78 ),
	.A(\UART_TX_Inst/n77 ));
   NAND2 \UART_TX_Inst/C225  (.OUT(\UART_TX_Inst/N139 ),
	.B(\UART_TX_Inst/n79 ),
	.A(\UART_TX_Inst/r31/AEQB [6]));
   NAND2 \UART_TX_Inst/C226  (.OUT(\UART_TX_Inst/N140 ),
	.B(\UART_TX_Inst/n80 ),
	.A(\UART_TX_Inst/r31/AEQB [5]));
   NAND2 \UART_TX_Inst/C227  (.OUT(\UART_TX_Inst/N141 ),
	.B(\UART_TX_Inst/n82 ),
	.A(\UART_TX_Inst/n81 ));
   NAND2 \UART_TX_Inst/C228  (.OUT(\UART_TX_Inst/N142 ),
	.B(\UART_TX_Inst/n84 ),
	.A(\UART_TX_Inst/n83 ));
   NAND2 \UART_TX_Inst/C229  (.OUT(\UART_TX_Inst/N143 ),
	.B(\UART_TX_Inst/n86 ),
	.A(\UART_TX_Inst/n85 ));
   NAND2 \UART_TX_Inst/C230  (.OUT(\UART_TX_Inst/N144 ),
	.B(\UART_TX_Inst/n87 ),
	.A(\UART_TX_Inst/r31/AEQB [1]));
   NAND2 \UART_TX_Inst/C231  (.OUT(\UART_TX_Inst/N145 ),
	.B(\UART_TX_Inst/n88 ),
	.A(\UART_TX_Inst/r_Clock_Count [0]));
   INV \UART_TX_Inst/I_6  (.OUT(\UART_TX_Inst/N146 ),
	.IN(\UART_TX_Inst/N145 ));
   INV \UART_TX_Inst/I_10  (.OUT(\UART_TX_Inst/N12 ),
	.IN(i_Rst_L));
   INV \UART_TX_Inst/I_13  (.OUT(\UART_TX_Inst/N18 ),
	.IN(\UART_TX_Inst/N17 ));
   NAND2 \UART_TX_Inst/lt_109/ULTI2  (.OUT(\UART_TX_Inst/N64 ),
	.B(\UART_TX_Inst/lt_109/LTV2 [2]),
	.A(\UART_TX_Inst/lt_109/LTV1 [2]));
   NAND2 \UART_TX_Inst/lt_109/ULTI1  (.OUT(\UART_TX_Inst/lt_109/LTV2 [2]),
	.B(\UART_TX_Inst/lt_109/LTV [2]),
	.A(\UART_TX_Inst/lt_109/AEQB [2]));
   NAND2 \UART_TX_Inst/lt_109/ULTI2_1  (.OUT(\UART_TX_Inst/lt_109/LTV [2]),
	.B(\UART_TX_Inst/lt_109/LTV2 [1]),
	.A(\UART_TX_Inst/lt_109/LTV1 [1]));
   NAND2 \UART_TX_Inst/lt_109/ULTI1_1  (.OUT(\UART_TX_Inst/lt_109/LTV2 [1]),
	.B(\UART_TX_Inst/lt_109/LTV [1]),
	.A(\UART_TX_Inst/lt_109/AEQB [1]));
   NAND2 \UART_TX_Inst/r31/ULTI1_1  (.OUT(\UART_TX_Inst/r31/LTV2 [1]),
	.B(\UART_TX_Inst/r31/LTV [1]),
	.A(\UART_TX_Inst/r31/AEQB [1]));
   NAND2 \UART_TX_Inst/r31/ULTI2_1  (.OUT(\UART_TX_Inst/r31/LTV [2]),
	.B(\UART_TX_Inst/r31/LTV2 [1]),
	.A(\UART_TX_Inst/r31/LTV1 [1]));
   NAND2 \UART_TX_Inst/r31/ULTI1_2  (.OUT(\UART_TX_Inst/r31/LTV2 [2]),
	.B(\UART_TX_Inst/r31/LTV [2]),
	.A(\UART_TX_Inst/r31/AEQB [2]));
   NAND2 \UART_TX_Inst/r31/ULTI1_3  (.OUT(\UART_TX_Inst/r31/LTV2 [3]),
	.B(\UART_TX_Inst/r31/LTV [3]),
	.A(\UART_TX_Inst/r31/AEQB [3]));
   NAND2 \UART_TX_Inst/r31/ULTI1_4  (.OUT(\UART_TX_Inst/r31/LTV2 [4]),
	.B(\UART_TX_Inst/r31/LTV [4]),
	.A(\UART_TX_Inst/r31/AEQB [4]));
   NAND2 \UART_TX_Inst/r31/ULTI1_5  (.OUT(\UART_TX_Inst/r31/LTV2 [5]),
	.B(\UART_TX_Inst/r31/LTV [5]),
	.A(\UART_TX_Inst/r31/AEQB [5]));
   NAND2 \UART_TX_Inst/r31/ULTI2_5  (.OUT(\UART_TX_Inst/r31/LTV [6]),
	.B(\UART_TX_Inst/r31/LTV2 [5]),
	.A(\UART_TX_Inst/r31/LTV1 [5]));
   NAND2 \UART_TX_Inst/r31/ULTI1_6  (.OUT(\UART_TX_Inst/r31/LTV2 [6]),
	.B(\UART_TX_Inst/r31/LTV [6]),
	.A(\UART_TX_Inst/r31/AEQB [6]));
   NAND2 \UART_TX_Inst/r31/ULTI2_6  (.OUT(\UART_TX_Inst/r31/LTV [7]),
	.B(\UART_TX_Inst/r31/LTV2 [6]),
	.A(\UART_TX_Inst/r31/LTV1 [6]));
   NAND2 \UART_TX_Inst/r31/ULTI1_7  (.OUT(\UART_TX_Inst/r31/LTV2 [7]),
	.B(\UART_TX_Inst/r31/LTV [7]),
	.A(\UART_TX_Inst/r31/AEQB [7]));
   NAND2 \UART_TX_Inst/r31/ULTI1_8  (.OUT(\UART_TX_Inst/r31/LTV2 [8]),
	.B(\UART_TX_Inst/r31/LTV [8]),
	.A(\UART_TX_Inst/r31/AEQB [8]));
   NAND2 \UART_TX_Inst/r31/ULTI2_8  (.OUT(\UART_TX_Inst/r31/LTV [9]),
	.B(\UART_TX_Inst/r31/LTV2 [8]),
	.A(\UART_TX_Inst/r31/LTV1 [8]));
   NAND2 \UART_TX_Inst/r31/ULTI1_9  (.OUT(\UART_TX_Inst/r31/LTV2 [9]),
	.B(\UART_TX_Inst/r31/LTV [9]),
	.A(\UART_TX_Inst/r31/AEQB [9]));
   NAND2 \UART_TX_Inst/r31/ULTI2_9  (.OUT(\UART_TX_Inst/r31/LTV [10]),
	.B(\UART_TX_Inst/r31/LTV2 [9]),
	.A(\UART_TX_Inst/r31/LTV1 [9]));
   NAND2 \UART_TX_Inst/r31/ULTI1  (.OUT(\UART_TX_Inst/r31/LTV2 [10]),
	.B(\UART_TX_Inst/r31/LTV [10]),
	.A(\UART_TX_Inst/r31/AEQB [10]));
   NAND2 \UART_RX_Inst/r35/ULTI0_0  (.OUT(\UART_RX_Inst/r35/LTV1 [0]),
	.B(\UART_RX_Inst/U3/U1/Z_9 ),
	.A(\UART_RX_Inst/N87 ));
   XNOR2 \UART_RX_Inst/r35/UEQI_1  (.OUT(\UART_RX_Inst/r35/AEQB [1]),
	.B(\UART_RX_Inst/U3/U1/Z_9 ),
	.A(\UART_RX_Inst/r_Clock_Count [1]));
   NAND2 \UART_RX_Inst/r35/ULTI0_1  (.OUT(\UART_RX_Inst/r35/LTV1 [1]),
	.B(\UART_RX_Inst/U3/U1/Z_9 ),
	.A(n71));
   NAND2 \UART_RX_Inst/r35/ULTI1_1  (.OUT(\UART_RX_Inst/r35/LTV2 [1]),
	.B(\UART_RX_Inst/r35/LTV [1]),
	.A(\UART_RX_Inst/r35/AEQB [1]));
   NAND2 \UART_RX_Inst/r35/ULTI2_1  (.OUT(\UART_RX_Inst/r35/LTV [2]),
	.B(\UART_RX_Inst/r35/LTV2 [1]),
	.A(\UART_RX_Inst/r35/LTV1 [1]));
   NAND2 \UART_RX_Inst/r35/ULTI1_2  (.OUT(\UART_RX_Inst/r35/LTV2 [2]),
	.B(\UART_RX_Inst/r35/LTV [2]),
	.A(\UART_RX_Inst/r35/AEQB [2]));
   NAND2 \UART_RX_Inst/r35/ULTI1_3  (.OUT(\UART_RX_Inst/r35/LTV2 [3]),
	.B(\UART_RX_Inst/r35/LTV [3]),
	.A(\UART_RX_Inst/r35/AEQB [3]));
   XNOR2 \UART_RX_Inst/r35/UEQI_4  (.OUT(\UART_RX_Inst/r35/AEQB [4]),
	.B(\UART_RX_Inst/U3/U1/Z_7 ),
	.A(\UART_RX_Inst/r_Clock_Count [4]));
   NAND2 \UART_RX_Inst/r35/ULTI0_4  (.OUT(\UART_RX_Inst/r35/LTV1 [4]),
	.B(\UART_RX_Inst/U3/U1/Z_7 ),
	.A(n68));
   NAND2 \UART_RX_Inst/r35/ULTI1_4  (.OUT(\UART_RX_Inst/r35/LTV2 [4]),
	.B(\UART_RX_Inst/r35/LTV [4]),
	.A(\UART_RX_Inst/r35/AEQB [4]));
   NAND2 \UART_RX_Inst/r35/ULTI2_4  (.OUT(\UART_RX_Inst/r35/LTV [5]),
	.B(\UART_RX_Inst/r35/LTV2 [4]),
	.A(\UART_RX_Inst/r35/LTV1 [4]));
   NAND2 \UART_RX_Inst/r35/ULTI1_5  (.OUT(\UART_RX_Inst/r35/LTV2 [5]),
	.B(\UART_RX_Inst/r35/LTV [5]),
	.A(\UART_RX_Inst/r35/AEQB [5]));
   NAND2 \UART_RX_Inst/r35/ULTI2_5  (.OUT(\UART_RX_Inst/r35/LTV [6]),
	.B(\UART_RX_Inst/r35/LTV2 [5]),
	.A(\UART_RX_Inst/r35/LTV1 [5]));
   XNOR2 \UART_RX_Inst/r35/UEQI_6  (.OUT(\UART_RX_Inst/r35/AEQB [6]),
	.B(\UART_RX_Inst/U3/U1/Z_9 ),
	.A(\UART_RX_Inst/r_Clock_Count [6]));
   NAND2 \UART_RX_Inst/r35/ULTI0_6  (.OUT(\UART_RX_Inst/r35/LTV1 [6]),
	.B(\UART_RX_Inst/U3/U1/Z_9 ),
	.A(n66));
   NAND2 \UART_RX_Inst/r35/ULTI1_6  (.OUT(\UART_RX_Inst/r35/LTV2 [6]),
	.B(\UART_RX_Inst/r35/LTV [6]),
	.A(\UART_RX_Inst/r35/AEQB [6]));
   NAND2 \UART_RX_Inst/r35/ULTI2_6  (.OUT(\UART_RX_Inst/r35/LTV [7]),
	.B(\UART_RX_Inst/r35/LTV2 [6]),
	.A(\UART_RX_Inst/r35/LTV1 [6]));
   XNOR2 \UART_RX_Inst/r35/UEQI_7  (.OUT(\UART_RX_Inst/r35/AEQB [7]),
	.B(\UART_RX_Inst/U3/U1/Z_7 ),
	.A(\UART_RX_Inst/r_Clock_Count [7]));
   NAND2 \UART_RX_Inst/r35/ULTI0_7  (.OUT(\UART_RX_Inst/r35/LTV1 [7]),
	.B(\UART_RX_Inst/U3/U1/Z_7 ),
	.A(n65));
   NAND2 \UART_RX_Inst/r35/ULTI1_7  (.OUT(\UART_RX_Inst/r35/LTV2 [7]),
	.B(\UART_RX_Inst/r35/LTV [7]),
	.A(\UART_RX_Inst/r35/AEQB [7]));
   NAND2 \UART_RX_Inst/r35/ULTI2_7  (.OUT(\UART_RX_Inst/r35/LTV [8]),
	.B(\UART_RX_Inst/r35/LTV2 [7]),
	.A(\UART_RX_Inst/r35/LTV1 [7]));
   NAND2 \UART_RX_Inst/r35/ULTI1_8  (.OUT(\UART_RX_Inst/r35/LTV2 [8]),
	.B(\UART_RX_Inst/r35/LTV [8]),
	.A(\UART_RX_Inst/r35/AEQB [8]));
   NAND2 \UART_RX_Inst/r35/ULTI2_8  (.OUT(\UART_RX_Inst/r35/LTV [9]),
	.B(\UART_RX_Inst/r35/LTV2 [8]),
	.A(\UART_RX_Inst/r35/LTV1 [8]));
   XNOR2 \UART_RX_Inst/r35/UEQI_9  (.OUT(\UART_RX_Inst/r35/AEQB [9]),
	.B(\UART_RX_Inst/U3/U1/Z_9 ),
	.A(\UART_RX_Inst/r_Clock_Count [9]));
   NAND2 \UART_RX_Inst/r35/ULTI0_9  (.OUT(\UART_RX_Inst/r35/LTV1 [9]),
	.B(\UART_RX_Inst/U3/U1/Z_9 ),
	.A(n63));
   NAND2 \UART_RX_Inst/r35/ULTI1_9  (.OUT(\UART_RX_Inst/r35/LTV2 [9]),
	.B(\UART_RX_Inst/r35/LTV [9]),
	.A(\UART_RX_Inst/r35/AEQB [9]));
   NAND2 \UART_RX_Inst/r35/ULTI2_9  (.OUT(\UART_RX_Inst/r35/LTV [10]),
	.B(\UART_RX_Inst/r35/LTV2 [9]),
	.A(\UART_RX_Inst/r35/LTV1 [9]));
   NAND2 \UART_RX_Inst/r35/ULTI1_10  (.OUT(\UART_RX_Inst/r35/LTV2 [10]),
	.B(\UART_RX_Inst/r35/LTV [10]),
	.A(\UART_RX_Inst/r35/AEQB [10]));
   NAND2 \UART_RX_Inst/r35/ULTI1_11  (.OUT(\UART_RX_Inst/r35/LTV2 [11]),
	.B(\UART_RX_Inst/r35/LTV [11]),
	.A(\UART_RX_Inst/r35/AEQB [11]));
   NAND2 \UART_RX_Inst/r35/ULTI1_12  (.OUT(\UART_RX_Inst/r35/LTV2 [12]),
	.B(\UART_RX_Inst/r35/LTV [12]),
	.A(\UART_RX_Inst/r35/AEQB [12]));
   NAND2 \UART_RX_Inst/r35/ULTI1_13  (.OUT(\UART_RX_Inst/r35/LTV2 [13]),
	.B(\UART_RX_Inst/r35/LTV [13]),
	.A(\UART_RX_Inst/r35/AEQB [13]));
   NAND2 \UART_RX_Inst/r35/ULTI1_14  (.OUT(\UART_RX_Inst/r35/LTV2 [14]),
	.B(\UART_RX_Inst/r35/LTV [14]),
	.A(\UART_RX_Inst/r35/AEQB [14]));
   NAND2 \UART_RX_Inst/r35/ULTI1  (.OUT(\UART_RX_Inst/r35/LTV2 [15]),
	.B(\UART_RX_Inst/r35/LTV [15]),
	.A(\UART_RX_Inst/r35/AEQB [15]));
   INV U1 (.OUT(\UART_TX_Inst/r31/LTV1 [0]),
	.IN(\UART_TX_Inst/N87 ));
   INV U2 (.OUT(\UART_TX_Inst/r31/LTV1 [1]),
	.IN(n80));
   INV U3 (.OUT(\UART_TX_Inst/r31/LTV1 [5]),
	.IN(n76));
   INV U4 (.OUT(\UART_TX_Inst/r31/LTV1 [6]),
	.IN(n75));
   INV U5 (.OUT(\UART_TX_Inst/r31/LTV1 [8]),
	.IN(n73));
   INV U6 (.OUT(\UART_TX_Inst/r31/LTV1 [9]),
	.IN(n72));
   INV U7 (.OUT(\UART_RX_Inst/r35/LTV1 [5]),
	.IN(n67));
   INV U8 (.OUT(\UART_RX_Inst/r35/LTV1 [8]),
	.IN(n64));
   INV U9 (.OUT(\UART_TX_Inst/r31/LTV [1]),
	.IN(\UART_TX_Inst/r31/LTV1 [0]));
   INV U10 (.OUT(\UART_TX_Inst/r31/LTV [3]),
	.IN(\UART_TX_Inst/r31/LTV2 [2]));
   INV U11 (.OUT(\UART_TX_Inst/r31/LTV [4]),
	.IN(\UART_TX_Inst/r31/LTV2 [3]));
   INV U12 (.OUT(\UART_TX_Inst/r31/LTV [5]),
	.IN(\UART_TX_Inst/r31/LTV2 [4]));
   INV U13 (.OUT(\UART_TX_Inst/r31/LTV [8]),
	.IN(\UART_TX_Inst/r31/LTV2 [7]));
   INV U14 (.OUT(\UART_TX_Inst/N23 ),
	.IN(\UART_TX_Inst/r31/LTV2 [10]));
   INV U15 (.OUT(\UART_RX_Inst/N145 ),
	.IN(\UART_RX_Inst/r35/LTV2 [15]));
   INV U16 (.OUT(\UART_RX_Inst/r35/LTV [1]),
	.IN(\UART_RX_Inst/r35/LTV1 [0]));
   INV U17 (.OUT(\UART_RX_Inst/r35/LTV [3]),
	.IN(\UART_RX_Inst/r35/LTV2 [2]));
   INV U18 (.OUT(\UART_RX_Inst/r35/LTV [4]),
	.IN(\UART_RX_Inst/r35/LTV2 [3]));
   INV U19 (.OUT(\UART_RX_Inst/r35/LTV [11]),
	.IN(\UART_RX_Inst/r35/LTV2 [10]));
   INV U20 (.OUT(\UART_RX_Inst/r35/LTV [12]),
	.IN(\UART_RX_Inst/r35/LTV2 [11]));
   INV U21 (.OUT(\UART_RX_Inst/r35/LTV [13]),
	.IN(\UART_RX_Inst/r35/LTV2 [12]));
   INV U22 (.OUT(\UART_RX_Inst/r35/LTV [14]),
	.IN(\UART_RX_Inst/r35/LTV2 [13]));
   INV U23 (.OUT(\UART_RX_Inst/r35/LTV [15]),
	.IN(\UART_RX_Inst/r35/LTV2 [14]));
   INV U24 (.OUT(\UART_TX_Inst/r31/AEQB [2]),
	.IN(\UART_TX_Inst/r_Clock_Count [2]));
   INV U25 (.OUT(\UART_TX_Inst/r31/AEQB [3]),
	.IN(\UART_TX_Inst/r_Clock_Count [3]));
   INV U26 (.OUT(\UART_TX_Inst/r31/AEQB [4]),
	.IN(\UART_TX_Inst/r_Clock_Count [4]));
   INV U27 (.OUT(\UART_TX_Inst/r31/AEQB [7]),
	.IN(\UART_TX_Inst/r_Clock_Count [7]));
   INV U28 (.OUT(\UART_TX_Inst/r31/AEQB [10]),
	.IN(\UART_TX_Inst/r_Clock_Count [10]));
   INV U29 (.OUT(\UART_RX_Inst/r35/AEQB [2]),
	.IN(\UART_RX_Inst/r_Clock_Count [2]));
   INV U30 (.OUT(\UART_RX_Inst/r35/AEQB [3]),
	.IN(\UART_RX_Inst/r_Clock_Count [3]));
   INV U31 (.OUT(\UART_RX_Inst/r35/AEQB [10]),
	.IN(\UART_RX_Inst/r_Clock_Count [10]));
   INV U32 (.OUT(\UART_RX_Inst/r35/AEQB [11]),
	.IN(\UART_RX_Inst/r_Clock_Count [11]));
   INV U33 (.OUT(\UART_RX_Inst/r35/AEQB [12]),
	.IN(\UART_RX_Inst/r_Clock_Count [12]));
   INV U34 (.OUT(\UART_RX_Inst/r35/AEQB [13]),
	.IN(\UART_RX_Inst/r_Clock_Count [13]));
   INV U35 (.OUT(\UART_RX_Inst/r35/AEQB [14]),
	.IN(\UART_RX_Inst/r_Clock_Count [14]));
   INV U36 (.OUT(\UART_RX_Inst/r35/AEQB [15]),
	.IN(\UART_RX_Inst/r_Clock_Count [15]));
   NOR2 U37 (.OUT(n1),
	.B(n2),
	.A(n74));
   NOR2 U38 (.OUT(n3),
	.B(n4),
	.A(n78));
   NOR2 U39 (.OUT(n5),
	.B(\UART_TX_Inst/N87 ),
	.A(n80));
   NOR2 U40 (.OUT(n6),
	.B(n7),
	.A(n61));
   NOR2 U41 (.OUT(n8),
	.B(n9),
	.A(n65));
   NOR2 U42 (.OUT(n10),
	.B(n11),
	.A(n69));
   NOR2 U43 (.OUT(n12),
	.B(\UART_RX_Inst/N87 ),
	.A(n71));
   NOR2 U44 (.OUT(n13),
	.B(n14),
	.A(n58));
   XNOR2 U45 (.OUT(n15),
	.B(n16),
	.A(\UART_TX_Inst/r_Clock_Count [10]));
   XNOR2 U46 (.OUT(n17),
	.B(n72),
	.A(n18));
   XNOR2 U47 (.OUT(\UART_TX_Inst/N95 ),
	.B(n1),
	.A(n73));
   XNOR2 U48 (.OUT(\UART_TX_Inst/N94 ),
	.B(n74),
	.A(n19));
   XNOR2 U49 (.OUT(\UART_TX_Inst/N93 ),
	.B(n21),
	.A(n20));
   XNOR2 U50 (.OUT(\UART_TX_Inst/N92 ),
	.B(n23),
	.A(n22));
   XNOR2 U51 (.OUT(\UART_TX_Inst/N91 ),
	.B(n3),
	.A(n77));
   XNOR2 U52 (.OUT(\UART_TX_Inst/N90 ),
	.B(n78),
	.A(n24));
   XNOR2 U53 (.OUT(\UART_TX_Inst/N89 ),
	.B(n5),
	.A(n79));
   XNOR2 U54 (.OUT(\UART_RX_Inst/N99 ),
	.B(n6),
	.A(n60));
   XNOR2 U55 (.OUT(\UART_RX_Inst/N98 ),
	.B(n61),
	.A(n25));
   XNOR2 U56 (.OUT(\UART_RX_Inst/N97 ),
	.B(n27),
	.A(n26));
   XNOR2 U57 (.OUT(\UART_RX_Inst/N96 ),
	.B(n29),
	.A(n28));
   XNOR2 U58 (.OUT(\UART_RX_Inst/N95 ),
	.B(n8),
	.A(n64));
   XNOR2 U59 (.OUT(\UART_RX_Inst/N94 ),
	.B(n65),
	.A(n30));
   XNOR2 U60 (.OUT(\UART_RX_Inst/N93 ),
	.B(n32),
	.A(n31));
   XNOR2 U61 (.OUT(\UART_RX_Inst/N92 ),
	.B(n34),
	.A(n33));
   XNOR2 U62 (.OUT(\UART_RX_Inst/N91 ),
	.B(n10),
	.A(n68));
   XNOR2 U63 (.OUT(\UART_RX_Inst/N90 ),
	.B(n69),
	.A(n35));
   XNOR2 U64 (.OUT(\UART_RX_Inst/N89 ),
	.B(n12),
	.A(n70));
   XNOR2 U65 (.OUT(\UART_RX_Inst/N102 ),
	.B(n13),
	.A(\UART_RX_Inst/n70 ));
   XNOR2 U66 (.OUT(\UART_RX_Inst/N101 ),
	.B(n36),
	.A(n58));
   XNOR2 U67 (.OUT(n37),
	.B(n59),
	.A(n38));
   NAND3 U68 (.OUT(n4),
	.C(n41),
	.B(n40),
	.A(n39));
   NAND3 U69 (.OUT(n22),
	.C(n24),
	.B(n43),
	.A(n42));
   NAND3 U70 (.OUT(n2),
	.C(n44),
	.B(n23),
	.A(n20));
   NAND3 U71 (.OUT(n18),
	.C(n19),
	.B(n46),
	.A(n45));
   NAND3 U72 (.OUT(n11),
	.C(n49),
	.B(n48),
	.A(n47));
   NAND3 U73 (.OUT(n33),
	.C(n35),
	.B(n51),
	.A(n50));
   NAND3 U74 (.OUT(n9),
	.C(n52),
	.B(n34),
	.A(n31));
   NAND3 U75 (.OUT(n28),
	.C(n30),
	.B(n54),
	.A(n53));
   NAND3 U76 (.OUT(n7),
	.C(n55),
	.B(n29),
	.A(n26));
   NAND3 U77 (.OUT(n38),
	.C(n25),
	.B(n57),
	.A(n56));
   NOR2 U78 (.OUT(n36),
	.B(n59),
	.A(n38));
   XNOR2 U79 (.OUT(\UART_TX_Inst/N88 ),
	.B(n40),
	.A(n80));
   XNOR2 U80 (.OUT(\UART_RX_Inst/N88 ),
	.B(n48),
	.A(n71));
   INV U81 (.OUT(n35),
	.IN(n11));
   INV U82 (.OUT(n52),
	.IN(n33));
   INV U83 (.OUT(n30),
	.IN(n9));
   INV U84 (.OUT(n55),
	.IN(n28));
   INV U85 (.OUT(n25),
	.IN(n7));
   INV U86 (.OUT(n24),
	.IN(n4));
   INV U87 (.OUT(n44),
	.IN(n22));
   INV U88 (.OUT(n19),
	.IN(n2));
   INV U89 (.OUT(n40),
	.IN(\UART_TX_Inst/N87 ));
   INV U90 (.OUT(n39),
	.IN(n80));
   INV U91 (.OUT(n41),
	.IN(n79));
   INV U92 (.OUT(n43),
	.IN(n78));
   INV U93 (.OUT(n42),
	.IN(n77));
   INV U94 (.OUT(n23),
	.IN(n76));
   INV U95 (.OUT(n20),
	.IN(n75));
   INV U96 (.OUT(n46),
	.IN(n74));
   INV U97 (.OUT(n45),
	.IN(n73));
   INV U98 (.OUT(n48),
	.IN(\UART_RX_Inst/N87 ));
   INV U99 (.OUT(n47),
	.IN(n71));
   INV U100 (.OUT(n49),
	.IN(n70));
   INV U101 (.OUT(n51),
	.IN(n69));
   INV U102 (.OUT(n50),
	.IN(n68));
   INV U103 (.OUT(n34),
	.IN(n67));
   INV U104 (.OUT(n31),
	.IN(n66));
   INV U105 (.OUT(n54),
	.IN(n65));
   INV U106 (.OUT(n53),
	.IN(n64));
   INV U107 (.OUT(n29),
	.IN(n63));
   INV U108 (.OUT(n26),
	.IN(n62));
   INV U109 (.OUT(n57),
	.IN(n61));
   INV U110 (.OUT(n56),
	.IN(n60));
   NOR2 U111 (.OUT(n16),
	.B(n72),
	.A(n18));
   NAND2 U112 (.OUT(n21),
	.B(n23),
	.A(n44));
   NAND2 U113 (.OUT(n27),
	.B(n29),
	.A(n55));
   NAND2 U114 (.OUT(n32),
	.B(n34),
	.A(n52));
   INV U115 (.OUT(n14),
	.IN(n36));
   INV U116 (.OUT(\UART_TX_Inst/N97 ),
	.IN(n15));
   INV U117 (.OUT(\UART_TX_Inst/N96 ),
	.IN(n17));
   INV U118 (.OUT(\UART_RX_Inst/N100 ),
	.IN(n37));
   INV U119 (.OUT(n58),
	.IN(\UART_RX_Inst/r_Clock_Count [14]));
   INV U120 (.OUT(n59),
	.IN(\UART_RX_Inst/r_Clock_Count [13]));
   INV U121 (.OUT(n60),
	.IN(\UART_RX_Inst/r_Clock_Count [12]));
   INV U122 (.OUT(n61),
	.IN(\UART_RX_Inst/r_Clock_Count [11]));
   INV U123 (.OUT(n62),
	.IN(\UART_RX_Inst/r_Clock_Count [10]));
   INV U124 (.OUT(n63),
	.IN(\UART_RX_Inst/r_Clock_Count [9]));
   INV U125 (.OUT(n64),
	.IN(\UART_RX_Inst/r35/AEQB [8]));
   INV U126 (.OUT(n65),
	.IN(\UART_RX_Inst/r_Clock_Count [7]));
   INV U127 (.OUT(n66),
	.IN(\UART_RX_Inst/r_Clock_Count [6]));
   INV U128 (.OUT(n67),
	.IN(\UART_RX_Inst/r35/AEQB [5]));
   INV U129 (.OUT(n68),
	.IN(\UART_RX_Inst/r_Clock_Count [4]));
   INV U130 (.OUT(n69),
	.IN(\UART_RX_Inst/r_Clock_Count [3]));
   INV U131 (.OUT(n70),
	.IN(\UART_RX_Inst/r_Clock_Count [2]));
   INV U132 (.OUT(n71),
	.IN(\UART_RX_Inst/r_Clock_Count [1]));
   INV U133 (.OUT(\UART_RX_Inst/N87 ),
	.IN(\UART_RX_Inst/r_Clock_Count [0]));
   INV U134 (.OUT(n72),
	.IN(\UART_TX_Inst/r31/AEQB [9]));
   INV U135 (.OUT(n73),
	.IN(\UART_TX_Inst/r31/AEQB [8]));
   INV U136 (.OUT(n74),
	.IN(\UART_TX_Inst/r_Clock_Count [7]));
   INV U137 (.OUT(n75),
	.IN(\UART_TX_Inst/r31/AEQB [6]));
   INV U138 (.OUT(n76),
	.IN(\UART_TX_Inst/r31/AEQB [5]));
   INV U139 (.OUT(n77),
	.IN(\UART_TX_Inst/r_Clock_Count [4]));
   INV U140 (.OUT(n78),
	.IN(\UART_TX_Inst/r_Clock_Count [3]));
   INV U141 (.OUT(n79),
	.IN(\UART_TX_Inst/r_Clock_Count [2]));
   INV U142 (.OUT(n80),
	.IN(\UART_TX_Inst/r31/AEQB [1]));
   INV U143 (.OUT(\UART_TX_Inst/N87 ),
	.IN(\UART_TX_Inst/r_Clock_Count [0]));
   INV U144 (.OUT(\UART_RX_Inst/lt_110/LTV1 [0]),
	.IN(\UART_RX_Inst/n168 ));
   INV U145 (.OUT(\UART_RX_Inst/lt_110/LTV1 [1]),
	.IN(\UART_RX_Inst/n167 ));
   INV U146 (.OUT(\UART_RX_Inst/lt_110/LTV1 [2]),
	.IN(\UART_RX_Inst/n166 ));
   INV U147 (.OUT(\UART_RX_Inst/lt_110/LTV [1]),
	.IN(\UART_RX_Inst/lt_110/LTV1 [0]));
   INV U148 (.OUT(\UART_TX_Inst/lt_109/LTV1 [0]),
	.IN(\UART_TX_Inst/N66 ));
   INV U149 (.OUT(\UART_TX_Inst/lt_109/LTV1 [1]),
	.IN(\UART_TX_Inst/n102 ));
   INV U150 (.OUT(\UART_TX_Inst/lt_109/LTV1 [2]),
	.IN(\UART_TX_Inst/n101 ));
   INV U151 (.OUT(\UART_TX_Inst/lt_109/LTV [1]),
	.IN(\UART_TX_Inst/lt_109/LTV1 [0]));
   INV U152 (.OUT(\UART_RX_Inst/n166 ),
	.IN(\UART_RX_Inst/lt_110/AEQB [2]));
   INV U153 (.OUT(\UART_TX_Inst/n101 ),
	.IN(\UART_TX_Inst/lt_109/AEQB [2]));
endmodule
