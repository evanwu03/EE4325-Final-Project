NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

DIVIDERCHAR "/" ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.042 ;
  SPACING 0.09 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M1

LAYER V1
  TYPE CUT ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M2

LAYER V2
  TYPE CUT ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M3

LAYER V3
  TYPE CUT ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M4

LAYER V4
  TYPE CUT ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M5

LAYER V5
  TYPE CUT ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
  END M6

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

SPACING
  SAMENET M1  M1    0.09 STACK ;
  SAMENET M2  M2    0.1 STACK ;
  SAMENET M3  M3    0.1 STACK ;
  SAMENET M4  M4    0.1 STACK ;
  SAMENET M5  M5    0.1 STACK ;
  SAMENET M6  M6    0.1 STACK ;
  SAMENET V1  V1    0.1 ;
  SAMENET V2  V2    0.1 ;
  SAMENET V3  V3    0.1 ;
  SAMENET V4  V4    0.1 ;
  SAMENET V5  V5    0.1 ;
  SAMENET V1  V2    0.00 STACK ;
  SAMENET V2  V3    0.00 STACK ;
  SAMENET V3  V4    0.00 STACK ;
  SAMENET V4  V5    0.00 STACK ;
  SAMENET V1  V3    0.00 STACK ;
  SAMENET V2  V4    0.00 STACK ;
  SAMENET V3  V5    0.00 STACK ;
  SAMENET V1  V4    0.00 STACK ;
  SAMENET V2  V5    0.00 STACK ;
  SAMENET V1  V5    0.00 STACK ;
END SPACING


VIA via5 DEFAULT
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5

VIA via4 DEFAULT
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4

VIA via3 DEFAULT
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3

VIA via2 DEFAULT
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2

VIA via1 DEFAULT
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1


VIARULE via1Array GENERATE
  LAYER M1 ;
  DIRECTION HORIZONTAL ;
  OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION VERTICAL ;
    OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER V1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via1Array


VIARULE via2Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via2Array


VIARULE via3Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER V5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via5Array

VIARULE TURNM1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
  LAYER M1 ;
    DIRECTION VERTICAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER M2 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER M3 ;
    DIRECTION VERTICAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE TURNM5 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
  LAYER M5 ;
    DIRECTION VERTICAL ;
END TURNM5

VIARULE TURNM6 GENERATE
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
END TURNM6


SITE  CoreSite
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.260 BY 5.98 ;
END  CoreSite

SITE  TDCoverSite
    CLASS       CORE ;
    SIZE        0.0500 BY 0.0500 ;
END  TDCoverSite

SITE  SBlockSite
    CLASS       CORE ;
    SIZE        0.0500 BY 0.0500 ;
END  SBlockSite

SITE  PortCellSite
    CLASS       PAD ;
    SIZE        0.0500 BY 0.0500 ;
END  PortCellSite

SITE  Core
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.260 BY 5.98 ;
END  Core



MACRO DFF
  CLASS CORE ;
  ORIGIN 4.427 2.002 ;
  FOREIGN DFF -4.427 -2.002 ;
  SIZE 8.32 BY 5.98 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -3.893 0.7 -3.751 1 ;
      LAYER M2 ;
        RECT -3.923 0.641 -3.702 1.027 ;
      LAYER V1 ;
        RECT -3.873 0.836 -3.773 0.936 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -2.022 0.7 -1.88 1 ;
      LAYER M2 ;
        RECT -2.032 0.641 -1.882 1.027 ;
      LAYER V1 ;
        RECT -2.004 0.836 -1.904 0.936 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.405 -0.957 3.515 2.805 ;
      LAYER M2 ;
        RECT 3.405 0.656 3.578 1.042 ;
      LAYER V1 ;
        RECT 3.409 0.851 3.509 0.951 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -3.086 0.7 -2.944 1 ;
      LAYER M2 ;
        RECT -3.072 0.641 -2.922 1.027 ;
      LAYER V1 ;
        RECT -3.064 0.836 -2.964 0.936 ;
    END
  END R
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -4.427 -2.002 3.893 -1.848 ;
        RECT 3.048 -2.002 3.158 -0.384 ;
        RECT 2.761 -2.002 2.871 -0.393 ;
        RECT 1.849 -2.002 1.959 -0.393 ;
        RECT 0.024 -2.002 0.134 -0.393 ;
        RECT -2.228 -2.002 -2.118 -0.393 ;
        RECT -3.081 -2.002 -2.971 -0.393 ;
        RECT -3.618 -2.002 -3.508 -0.379 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -4.427 3.835 3.893 3.978 ;
        RECT 3.037 1.82 3.147 3.978 ;
        RECT 1.828 1.832 1.938 3.978 ;
        RECT 0.003 1.832 0.113 3.978 ;
        RECT -2.133 1.832 -2.023 3.978 ;
        RECT -3.618 1.832 -3.508 3.978 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 2.753 1.409 2.863 2.798 ;
      RECT 1.608 1.409 2.863 1.519 ;
      RECT 1.2 1.182 2.712 1.292 ;
      RECT 1.2 0.961 1.31 1.292 ;
      RECT -1.522 0.961 1.31 1.071 ;
      RECT -1.522 0.485 -1.412 1.071 ;
      RECT -2.958 0.485 -1.412 0.595 ;
      RECT -0.792 0.582 2.487 0.692 ;
      RECT 2.377 -0.095 2.487 0.692 ;
      RECT 1.327 -0.095 2.487 0.015 ;
      RECT 1.622 -0.3 2.455 -0.19 ;
      RECT 2.345 -0.95 2.455 -0.19 ;
      RECT 1.014 1.627 1.124 2.812 ;
      RECT 1.014 1.627 2.239 1.737 ;
      RECT 1.045 0.258 2.236 0.368 ;
      RECT 1.045 -0.952 1.155 0.368 ;
      RECT -3.348 -0.957 -3.238 2.797 ;
      RECT -3.348 0.265 0.861 0.375 ;
      RECT -1.228 3.009 -0.403 3.119 ;
      RECT -0.513 1.426 -0.403 3.119 ;
      RECT -0.513 1.426 0.861 1.536 ;
      RECT -3.089 1.217 -2.979 2.802 ;
      RECT -3.089 1.217 -0.179 1.327 ;
      RECT -2.705 -0.033 -0.194 0.077 ;
      RECT -2.705 -0.956 -2.595 0.077 ;
      RECT -1.43 3.245 -0.707 3.355 ;
      RECT -1.43 1.617 -1.32 3.355 ;
      RECT -3.411 2.95 -2.402 3.06 ;
      RECT -2.512 1.617 -2.402 3.06 ;
      RECT -2.512 1.617 -1.32 1.727 ;
      RECT -2.358 -0.234 -0.948 -0.124 ;
      RECT -1.058 -0.95 -0.948 -0.124 ;
      RECT -1.086 1.417 -0.976 2.804 ;
      RECT -2.338 1.417 -0.976 1.527 ;
      RECT -4.128 -0.957 -4.018 2.797 ;
      RECT -4.128 0.428 -3.455 0.538 ;
      RECT 2.152 0.866 3.228 0.976 ;
  END
 
END DFF

MACRO FILLER
  CLASS CORE ;
  ORIGIN 0.263 3.998 ;
  FOREIGN FILLER -0.263 -3.998 ;
  SIZE 0.26 BY 5.98 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.363 -3.998 0.097 -3.844 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.363 1.839 0.097 1.982 ;
    END
  END VDD!
 
END FILLER

MACRO INV
  CLASS CORE ;
  ORIGIN 0.618 2.538 ;
  FOREIGN INV -0.618 -2.538 ;
  SIZE 1.3 BY 5.98 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.3 0.128 -0.158 0.428 ;
      LAYER M2 ;
        RECT -0.303 0.12 -0.153 0.506 ;
      LAYER V1 ;
        RECT -0.28 0.264 -0.18 0.364 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 -1.498 0.352 2.257 ;
      LAYER M2 ;
        RECT 0.217 0.12 0.367 0.506 ;
      LAYER V1 ;
        RECT 0.25 0.264 0.35 0.364 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.618 -2.538 0.682 -2.384 ;
        RECT -0.311 -2.538 -0.201 -0.925 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.618 3.299 0.682 3.442 ;
        RECT -0.305 1.295 -0.195 3.442 ;
    END
  END VDD!
  
END INV

MACRO NAND2
  CLASS CORE ;
  ORIGIN 0.916 2.835 ;
  FOREIGN NAND2 -0.916 -2.835 ;
  SIZE 2.08 BY 5.98 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.337 -0.172 -0.195 0.128 ;
      LAYER M2 ;
        RECT -0.341 -0.177 -0.191 0.209 ;
      LAYER V1 ;
        RECT -0.315 -0.036 -0.215 0.064 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.183 -0.17 0.325 0.13 ;
      LAYER M2 ;
        RECT 0.179 -0.177 0.329 0.209 ;
      LAYER V1 ;
        RECT 0.206 -0.034 0.306 0.066 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.736 -0.112 0.846 1.96 ;
        RECT -0.625 0.583 0.846 0.693 ;
        RECT -0.625 -1.785 -0.515 1.96 ;
      LAYER M2 ;
        RECT 0.699 -0.177 0.849 0.209 ;
      LAYER V1 ;
        RECT 0.742 -0.067 0.842 0.033 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.916 -2.835 1.164 -2.681 ;
        RECT 0.728 -2.835 0.838 -1.228 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.916 3.002 1.164 3.145 ;
        RECT -0.232 1.004 -0.122 3.145 ;
    END
  END VDD!
  
END NAND2

MACRO NAND3
  CLASS CORE ;
  ORIGIN 1.273 2.268 ;
  FOREIGN NAND3 -1.273 -2.268 ;
  SIZE 2.6 BY 5.98 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.693 0.4 -0.551 0.7 ;
      LAYER M2 ;
        RECT -0.698 0.39 -0.548 0.776 ;
      LAYER V1 ;
        RECT -0.671 0.536 -0.571 0.636 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.174 0.393 -0.032 0.693 ;
      LAYER M2 ;
        RECT -0.178 0.39 -0.028 0.776 ;
      LAYER V1 ;
        RECT -0.152 0.529 -0.052 0.629 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.867 0.402 1.009 0.702 ;
      LAYER M2 ;
        RECT 0.862 0.39 1.012 0.776 ;
      LAYER V1 ;
        RECT 0.889 0.538 0.989 0.638 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.901 0.971 1.011 2.536 ;
        RECT -0.964 0.971 1.011 1.081 ;
        RECT 0.376 0.399 0.486 1.081 ;
        RECT -0.571 0.971 -0.461 2.532 ;
        RECT -0.964 -1.218 -0.854 1.081 ;
      LAYER M2 ;
        RECT 0.342 0.39 0.492 0.776 ;
      LAYER V1 ;
        RECT 0.378 0.527 0.478 0.627 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -1.273 -2.268 1.327 -2.114 ;
        RECT 0.907 -2.268 1.017 -0.646 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -1.273 3.569 1.327 3.712 ;
        RECT 0.41 1.569 0.52 3.712 ;
        RECT -0.964 1.565 -0.854 3.712 ;
    END
  END VDD!
 
END NAND3

MACRO NOR2
  CLASS CORE ;
  ORIGIN 1.149 2.627 ;
  FOREIGN NOR2 -1.149 -2.627 ;
  SIZE 2.08 BY 5.98 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.57 0.043 -0.428 0.343 ;
      LAYER M2 ;
        RECT -0.574 0.031 -0.424 0.417 ;
      LAYER V1 ;
        RECT -0.548 0.179 -0.448 0.279 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.05 0.043 0.092 0.343 ;
      LAYER M2 ;
        RECT -0.054 0.031 0.096 0.417 ;
      LAYER V1 ;
        RECT -0.027 0.179 0.073 0.279 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.508 -0.272 0.618 2.17 ;
        RECT -0.295 -0.272 0.618 -0.162 ;
        RECT -0.295 -1.584 -0.185 -0.162 ;
      LAYER M2 ;
        RECT 0.466 0.031 0.616 0.417 ;
      LAYER V1 ;
        RECT 0.509 0.179 0.609 0.279 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -1.149 -2.627 0.931 -2.473 ;
        RECT 0.497 -2.627 0.607 -1.021 ;
        RECT -0.858 -2.627 -0.748 -1.01 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -1.149 3.21 0.931 3.353 ;
        RECT -0.858 1.208 -0.748 3.353 ;
    END
  END VDD!
  
END NOR2

MACRO OAI22
  CLASS CORE ;
  ORIGIN 1.401 1.167 ;
  FOREIGN OAI22 -1.401 -1.167 ;
  SIZE 2.86 BY 5.98 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -1.101 1.5 -0.959 1.8 ;
      LAYER M2 ;
        RECT -1.086 1.491 -0.936 1.877 ;
      LAYER V1 ;
        RECT -1.079 1.636 -0.979 1.736 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.564 1.5 -0.422 1.8 ;
      LAYER M2 ;
        RECT -0.566 1.491 -0.416 1.877 ;
      LAYER V1 ;
        RECT -0.541 1.636 -0.441 1.736 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.996 1.5 1.138 1.8 ;
      LAYER M2 ;
        RECT 0.994 1.491 1.144 1.877 ;
      LAYER V1 ;
        RECT 1.02 1.636 1.12 1.736 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.044 1.5 0.098 1.8 ;
      LAYER M2 ;
        RECT -0.046 1.491 0.104 1.877 ;
      LAYER V1 ;
        RECT -0.02 1.636 0.08 1.736 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.494 1.493 0.604 2.134 ;
        RECT -0.136 2.024 0.604 2.134 ;
        RECT -0.136 2.024 -0.026 3.621 ;
        RECT -0.827 2.025 -0.026 2.135 ;
        RECT -0.827 -0.207 -0.717 2.135 ;
      LAYER M2 ;
        RECT 0.474 1.491 0.624 1.877 ;
      LAYER V1 ;
        RECT 0.5 1.631 0.6 1.731 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -1.401 -1.167 1.459 -1.013 ;
        RECT 0.437 -1.167 0.547 0.437 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -1.401 4.67 1.459 4.813 ;
        RECT 0.988 2.666 1.098 4.813 ;
        RECT -1.092 2.668 -0.982 4.813 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT -0.146 0.604 1.011 0.714 ;
      RECT 0.901 -0.118 1.011 0.714 ;
      RECT -0.146 -0.507 -0.036 0.714 ;
      RECT -1.097 -0.507 -0.987 0.444 ;
      RECT -1.097 -0.507 -0.036 -0.397 ;
  END
  
END OAI22

MACRO XNOR2
  CLASS CORE ;
  ORIGIN 1.21 0.964 ;
  FOREIGN XNOR2 -1.21 -0.964 ;
  SIZE 2.86 BY 5.98 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.197 1.702 1.339 2.002 ;
      LAYER M2 ;
        RECT 1.185 1.694 1.335 2.08 ;
      LAYER V1 ;
        RECT 1.213 1.865 1.313 1.965 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.366 1.728 -0.224 2.028 ;
      LAYER M2 ;
        RECT -0.375 1.694 -0.225 2.08 ;
      LAYER V1 ;
        RECT -0.344 1.864 -0.244 1.964 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.433 0.728 1.049 0.838 ;
        RECT 0.939 0.095 1.049 0.838 ;
        RECT 0.433 0.728 0.543 3.83 ;
      LAYER M2 ;
        RECT 0.405 1.694 0.555 2.08 ;
      LAYER V1 ;
        RECT 0.438 1.848 0.538 1.948 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -1.21 -0.964 1.65 -0.81 ;
        RECT -0.104 -0.964 0.006 0.645 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -1.21 4.873 1.65 5.016 ;
        RECT 1.205 2.872 1.315 5.016 ;
        RECT -0.092 2.872 0.018 5.016 ;
        RECT -0.935 2.875 -0.825 5.016 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.207 -0.204 1.317 0.644 ;
      RECT 0.425 -0.204 0.535 0.637 ;
      RECT 0.425 -0.204 1.317 -0.094 ;
      RECT -0.647 2.254 -0.537 3.841 ;
      RECT -0.935 2.254 0.254 2.364 ;
      RECT -0.935 0.086 -0.825 2.364 ;
  END
  
END XNOR2

END LIBRARY
