module inv(in, out);
input in;
output out;
//assign out = ~in;
endmodule

module nand2(a, b, out);
input a, b;
output out;
// out = ~(a & b);
endmodule

module nand3(a, b, c, out);
input a, b, c;
output out;
//assign out = ~(a & b & c);
endmodule

module nand4(a, b, c, d, out);
input a, b, c, d;
output out;
//assign out = ~(a & b & c & d);
endmodule

module nor2(a, b, out);
input a, b;
output out;
//assign out = ~(a | b);
endmodule

module nor3(a, b, c, out);
input a, b, c;
output out;
//assign out = ~(a | b | c);
endmodule

module xor2(a, b, out);
input a, b;
output out;
//assign out = (a ^ b);
endmodule

module aoi12(a, b, c, out);
input a, b, c;
output out;
//assign out = ~(a | (b & c));
endmodule

module aoi22(a, b, c, d, out);
input a, b, c, d;
output out;
//assign out = ~((a & b) | (c & d));
endmodule

module oai12(a, b, c, out);
input a, b, c;
output out;
//assign out = ~(a & (b | c));
endmodule

module oai22(a, b, c, d, out);
input a, b, c, d;
output out;
//assign out = ~((a | b) & (c | d));
endmodule

module dff( d, gclk, rnot, q);
input d, gclk, rnot;
output q;
reg q;
/*
always @(posedge gclk or negedge rnot)
  if (rnot == 1'b0)
    q = 1'b0;
  else
    q = d;
*/
endmodule


