* File: inv.pex.sp
* Created: Mon Apr 14 11:47:27 2025
* Program "Calibre xRC"
* Version "v2024.4_12.9"
* 
.include "inv.pex.sp.pex"
.subckt inv  GND! OUT VDD! INA
* 
* INA	INA
* VDD!	VDD!
* OUT	OUT
* GND!	GND!
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=3.5464e-12
+ PERIM=8.056e-06
XMMN0 N_OUT_MMN0_d N_INA_MMN0_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET
+ L=6.5e-08 W=5.6e-07 AD=2.1616e-13 AS=1.232e-13 PD=1.892e-06 PS=1.56e-06
+ NRD=0.576786 NRS=0.283929 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=2.2e-07 SB=3.86e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=1.1505e-14 PANW9=2.4895e-14 PANW10=0
XMMP0 N_OUT_MMP0_d N_INA_MMP0_g N_VDD!_MMP0_s N_VDD!_D0_noxref_neg PFET
+ L=6.5e-08 W=9.55e-07 AD=3.6863e-13 AS=2.101e-13 PD=2.682e-06 PS=2.35e-06
+ NRD=0.33822 NRS=0.164398 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=2.2e-07 SB=3.86e-07 SD=0 PANW1=4.615e-15 PANW2=3.25e-15 PANW3=3.25e-15
+ PANW4=3.25e-15 PANW5=3.25e-15 PANW6=6.8575e-14 PANW7=7.5075e-14 PANW8=1.3e-14
+ PANW9=1.196e-14 PANW10=2.964e-14
*
.include "inv.pex.sp.INV.pxi"
*
.ends
*
*
